magic
tech sky130A
magscale 1 2
timestamp 1730624594
<< pwell >>
rect -246 -737 246 737
<< nmos >>
rect -50 427 50 527
rect -50 109 50 209
rect -50 -209 50 -109
rect -50 -527 50 -427
<< ndiff >>
rect -108 515 -50 527
rect -108 439 -96 515
rect -62 439 -50 515
rect -108 427 -50 439
rect 50 515 108 527
rect 50 439 62 515
rect 96 439 108 515
rect 50 427 108 439
rect -108 197 -50 209
rect -108 121 -96 197
rect -62 121 -50 197
rect -108 109 -50 121
rect 50 197 108 209
rect 50 121 62 197
rect 96 121 108 197
rect 50 109 108 121
rect -108 -121 -50 -109
rect -108 -197 -96 -121
rect -62 -197 -50 -121
rect -108 -209 -50 -197
rect 50 -121 108 -109
rect 50 -197 62 -121
rect 96 -197 108 -121
rect 50 -209 108 -197
rect -108 -439 -50 -427
rect -108 -515 -96 -439
rect -62 -515 -50 -439
rect -108 -527 -50 -515
rect 50 -439 108 -427
rect 50 -515 62 -439
rect 96 -515 108 -439
rect 50 -527 108 -515
<< ndiffc >>
rect -96 439 -62 515
rect 62 439 96 515
rect -96 121 -62 197
rect 62 121 96 197
rect -96 -197 -62 -121
rect 62 -197 96 -121
rect -96 -515 -62 -439
rect 62 -515 96 -439
<< psubdiff >>
rect -210 667 -114 701
rect 114 667 210 701
rect -210 605 -176 667
rect 176 605 210 667
rect -210 -667 -176 -605
rect 176 -667 210 -605
rect -210 -701 -114 -667
rect 114 -701 210 -667
<< psubdiffcont >>
rect -114 667 114 701
rect -210 -605 -176 605
rect 176 -605 210 605
rect -114 -701 114 -667
<< poly >>
rect -50 599 50 615
rect -50 565 -34 599
rect 34 565 50 599
rect -50 527 50 565
rect -50 389 50 427
rect -50 355 -34 389
rect 34 355 50 389
rect -50 339 50 355
rect -50 281 50 297
rect -50 247 -34 281
rect 34 247 50 281
rect -50 209 50 247
rect -50 71 50 109
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -109 50 -71
rect -50 -247 50 -209
rect -50 -281 -34 -247
rect 34 -281 50 -247
rect -50 -297 50 -281
rect -50 -355 50 -339
rect -50 -389 -34 -355
rect 34 -389 50 -355
rect -50 -427 50 -389
rect -50 -565 50 -527
rect -50 -599 -34 -565
rect 34 -599 50 -565
rect -50 -615 50 -599
<< polycont >>
rect -34 565 34 599
rect -34 355 34 389
rect -34 247 34 281
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -281 34 -247
rect -34 -389 34 -355
rect -34 -599 34 -565
<< locali >>
rect -210 667 -114 701
rect 114 667 210 701
rect -210 605 -176 667
rect 176 605 210 667
rect -50 565 -34 599
rect 34 565 50 599
rect -96 515 -62 531
rect -96 423 -62 439
rect 62 515 96 531
rect 62 423 96 439
rect -50 355 -34 389
rect 34 355 50 389
rect -50 247 -34 281
rect 34 247 50 281
rect -96 197 -62 213
rect -96 105 -62 121
rect 62 197 96 213
rect 62 105 96 121
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -121 -62 -105
rect -96 -213 -62 -197
rect 62 -121 96 -105
rect 62 -213 96 -197
rect -50 -281 -34 -247
rect 34 -281 50 -247
rect -50 -389 -34 -355
rect 34 -389 50 -355
rect -96 -439 -62 -423
rect -96 -531 -62 -515
rect 62 -439 96 -423
rect 62 -531 96 -515
rect -50 -599 -34 -565
rect 34 -599 50 -565
rect -210 -667 -176 -605
rect 176 -667 210 -605
rect -210 -701 -114 -667
rect 114 -701 210 -667
<< viali >>
rect -34 565 34 599
rect -96 439 -62 515
rect 62 439 96 515
rect -34 355 34 389
rect -34 247 34 281
rect -96 121 -62 197
rect 62 121 96 197
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -197 -62 -121
rect 62 -197 96 -121
rect -34 -281 34 -247
rect -34 -389 34 -355
rect -96 -515 -62 -439
rect 62 -515 96 -439
rect -34 -599 34 -565
<< metal1 >>
rect -46 599 46 605
rect -46 565 -34 599
rect 34 565 46 599
rect -46 559 46 565
rect -102 515 -56 527
rect -102 439 -96 515
rect -62 439 -56 515
rect -102 427 -56 439
rect 56 515 102 527
rect 56 439 62 515
rect 96 439 102 515
rect 56 427 102 439
rect -46 389 46 395
rect -46 355 -34 389
rect 34 355 46 389
rect -46 349 46 355
rect -46 281 46 287
rect -46 247 -34 281
rect 34 247 46 281
rect -46 241 46 247
rect -102 197 -56 209
rect -102 121 -96 197
rect -62 121 -56 197
rect -102 109 -56 121
rect 56 197 102 209
rect 56 121 62 197
rect 96 121 102 197
rect 56 109 102 121
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -121 -56 -109
rect -102 -197 -96 -121
rect -62 -197 -56 -121
rect -102 -209 -56 -197
rect 56 -121 102 -109
rect 56 -197 62 -121
rect 96 -197 102 -121
rect 56 -209 102 -197
rect -46 -247 46 -241
rect -46 -281 -34 -247
rect 34 -281 46 -247
rect -46 -287 46 -281
rect -46 -355 46 -349
rect -46 -389 -34 -355
rect 34 -389 46 -355
rect -46 -395 46 -389
rect -102 -439 -56 -427
rect -102 -515 -96 -439
rect -62 -515 -56 -439
rect -102 -527 -56 -515
rect 56 -439 102 -427
rect 56 -515 62 -439
rect 96 -515 102 -439
rect 56 -527 102 -515
rect -46 -565 46 -559
rect -46 -599 -34 -565
rect 34 -599 46 -565
rect -46 -605 46 -599
<< properties >>
string FIXED_BBOX -193 -684 193 684
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.5 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
