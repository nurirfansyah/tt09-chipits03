magic
tech sky130A
magscale 1 2
timestamp 1730448391
<< error_p >>
rect -29 635 29 641
rect -29 601 -17 635
rect -29 595 29 601
rect -29 407 29 413
rect -29 373 -17 407
rect -29 367 29 373
rect -29 299 29 305
rect -29 265 -17 299
rect -29 259 29 265
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -265 29 -259
rect -29 -299 -17 -265
rect -29 -305 29 -299
rect -29 -373 29 -367
rect -29 -407 -17 -373
rect -29 -413 29 -407
rect -29 -601 29 -595
rect -29 -635 -17 -601
rect -29 -641 29 -635
<< nwell >>
rect -211 -773 211 773
<< pmos >>
rect -15 454 15 554
rect -15 118 15 218
rect -15 -218 15 -118
rect -15 -554 15 -454
<< pdiff >>
rect -73 542 -15 554
rect -73 466 -61 542
rect -27 466 -15 542
rect -73 454 -15 466
rect 15 542 73 554
rect 15 466 27 542
rect 61 466 73 542
rect 15 454 73 466
rect -73 206 -15 218
rect -73 130 -61 206
rect -27 130 -15 206
rect -73 118 -15 130
rect 15 206 73 218
rect 15 130 27 206
rect 61 130 73 206
rect 15 118 73 130
rect -73 -130 -15 -118
rect -73 -206 -61 -130
rect -27 -206 -15 -130
rect -73 -218 -15 -206
rect 15 -130 73 -118
rect 15 -206 27 -130
rect 61 -206 73 -130
rect 15 -218 73 -206
rect -73 -466 -15 -454
rect -73 -542 -61 -466
rect -27 -542 -15 -466
rect -73 -554 -15 -542
rect 15 -466 73 -454
rect 15 -542 27 -466
rect 61 -542 73 -466
rect 15 -554 73 -542
<< pdiffc >>
rect -61 466 -27 542
rect 27 466 61 542
rect -61 130 -27 206
rect 27 130 61 206
rect -61 -206 -27 -130
rect 27 -206 61 -130
rect -61 -542 -27 -466
rect 27 -542 61 -466
<< nsubdiff >>
rect -175 703 -79 737
rect 79 703 175 737
rect -175 641 -141 703
rect 141 641 175 703
rect -175 -703 -141 -641
rect 141 -703 175 -641
rect -175 -737 -79 -703
rect 79 -737 175 -703
<< nsubdiffcont >>
rect -79 703 79 737
rect -175 -641 -141 641
rect 141 -641 175 641
rect -79 -737 79 -703
<< poly >>
rect -33 635 33 651
rect -33 601 -17 635
rect 17 601 33 635
rect -33 585 33 601
rect -15 554 15 585
rect -15 423 15 454
rect -33 407 33 423
rect -33 373 -17 407
rect 17 373 33 407
rect -33 357 33 373
rect -33 299 33 315
rect -33 265 -17 299
rect 17 265 33 299
rect -33 249 33 265
rect -15 218 15 249
rect -15 87 15 118
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -118 15 -87
rect -15 -249 15 -218
rect -33 -265 33 -249
rect -33 -299 -17 -265
rect 17 -299 33 -265
rect -33 -315 33 -299
rect -33 -373 33 -357
rect -33 -407 -17 -373
rect 17 -407 33 -373
rect -33 -423 33 -407
rect -15 -454 15 -423
rect -15 -585 15 -554
rect -33 -601 33 -585
rect -33 -635 -17 -601
rect 17 -635 33 -601
rect -33 -651 33 -635
<< polycont >>
rect -17 601 17 635
rect -17 373 17 407
rect -17 265 17 299
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -299 17 -265
rect -17 -407 17 -373
rect -17 -635 17 -601
<< locali >>
rect -175 703 -79 737
rect 79 703 175 737
rect -175 641 -141 703
rect 141 641 175 703
rect -33 601 -17 635
rect 17 601 33 635
rect -61 542 -27 558
rect -61 450 -27 466
rect 27 542 61 558
rect 27 450 61 466
rect -33 373 -17 407
rect 17 373 33 407
rect -33 265 -17 299
rect 17 265 33 299
rect -61 206 -27 222
rect -61 114 -27 130
rect 27 206 61 222
rect 27 114 61 130
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -130 -27 -114
rect -61 -222 -27 -206
rect 27 -130 61 -114
rect 27 -222 61 -206
rect -33 -299 -17 -265
rect 17 -299 33 -265
rect -33 -407 -17 -373
rect 17 -407 33 -373
rect -61 -466 -27 -450
rect -61 -558 -27 -542
rect 27 -466 61 -450
rect 27 -558 61 -542
rect -33 -635 -17 -601
rect 17 -635 33 -601
rect -175 -703 -141 -641
rect 141 -703 175 -641
rect -175 -737 -79 -703
rect 79 -737 175 -703
<< viali >>
rect -17 601 17 635
rect -61 466 -27 542
rect 27 466 61 542
rect -17 373 17 407
rect -17 265 17 299
rect -61 130 -27 206
rect 27 130 61 206
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -206 -27 -130
rect 27 -206 61 -130
rect -17 -299 17 -265
rect -17 -407 17 -373
rect -61 -542 -27 -466
rect 27 -542 61 -466
rect -17 -635 17 -601
<< metal1 >>
rect -29 635 29 641
rect -29 601 -17 635
rect 17 601 29 635
rect -29 595 29 601
rect -67 542 -21 554
rect -67 466 -61 542
rect -27 466 -21 542
rect -67 454 -21 466
rect 21 542 67 554
rect 21 466 27 542
rect 61 466 67 542
rect 21 454 67 466
rect -29 407 29 413
rect -29 373 -17 407
rect 17 373 29 407
rect -29 367 29 373
rect -29 299 29 305
rect -29 265 -17 299
rect 17 265 29 299
rect -29 259 29 265
rect -67 206 -21 218
rect -67 130 -61 206
rect -27 130 -21 206
rect -67 118 -21 130
rect 21 206 67 218
rect 21 130 27 206
rect 61 130 67 206
rect 21 118 67 130
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -130 -21 -118
rect -67 -206 -61 -130
rect -27 -206 -21 -130
rect -67 -218 -21 -206
rect 21 -130 67 -118
rect 21 -206 27 -130
rect 61 -206 67 -130
rect 21 -218 67 -206
rect -29 -265 29 -259
rect -29 -299 -17 -265
rect 17 -299 29 -265
rect -29 -305 29 -299
rect -29 -373 29 -367
rect -29 -407 -17 -373
rect 17 -407 29 -373
rect -29 -413 29 -407
rect -67 -466 -21 -454
rect -67 -542 -61 -466
rect -27 -542 -21 -466
rect -67 -554 -21 -542
rect 21 -466 67 -454
rect 21 -542 27 -466
rect 61 -542 67 -466
rect 21 -554 67 -542
rect -29 -601 29 -595
rect -29 -635 -17 -601
rect 17 -635 29 -601
rect -29 -641 29 -635
<< properties >>
string FIXED_BBOX -158 -720 158 720
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.5 l 0.15 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
