magic
tech sky130A
magscale 1 2
timestamp 1729033186
<< error_s >>
rect 126 628 284 637
rect 126 603 343 628
rect 55 123 64 603
rect 89 517 118 603
rect 185 594 343 603
rect 89 225 123 517
rect 209 505 222 535
rect 238 526 265 535
rect 247 505 260 526
rect 363 508 475 638
rect 917 628 1075 637
rect 917 603 1134 628
rect 207 501 234 505
rect 235 501 262 505
rect 207 495 297 501
rect 231 492 297 495
rect 235 491 262 492
rect 235 486 293 491
rect 231 476 262 485
rect 249 467 262 476
rect 144 463 157 467
rect 169 463 178 467
rect 232 463 266 467
rect 132 263 178 463
rect 220 461 278 463
rect 226 458 278 461
rect 203 453 212 458
rect 234 454 278 458
rect 291 454 300 458
rect 192 442 220 453
rect 234 451 272 454
rect 232 442 272 451
rect 203 275 272 442
rect 285 442 300 454
rect 312 454 325 458
rect 203 266 237 275
rect 203 263 212 266
rect 220 263 235 266
rect 249 263 279 275
rect 144 259 157 263
rect 169 259 178 263
rect 191 259 279 263
rect 148 254 279 259
rect 285 266 304 442
rect 285 254 300 266
rect 203 250 237 254
rect 176 225 234 231
rect 249 228 279 254
rect 291 250 300 254
rect 312 254 337 454
rect 346 254 475 508
rect 545 500 603 506
rect 545 466 557 500
rect 545 460 603 466
rect 312 250 325 254
rect 89 177 118 225
rect 172 216 238 225
rect 346 216 359 254
rect 176 210 188 216
rect 363 210 475 254
rect 172 191 238 210
rect 176 185 234 191
rect 346 185 475 210
rect 89 176 123 177
rect 89 142 346 176
rect 55 108 346 123
rect 363 106 475 185
rect 545 172 603 178
rect 545 138 557 172
rect 545 132 603 138
rect 846 123 855 603
rect 880 517 909 603
rect 976 594 1134 603
rect 880 225 914 517
rect 1000 505 1013 535
rect 1029 526 1056 535
rect 1038 505 1051 526
rect 1154 508 1266 638
rect 1708 628 1866 637
rect 1708 603 1925 628
rect 998 501 1025 505
rect 1026 501 1053 505
rect 998 495 1088 501
rect 1022 492 1088 495
rect 1026 491 1053 492
rect 1026 486 1084 491
rect 1022 476 1053 485
rect 1040 467 1053 476
rect 935 463 948 467
rect 960 463 969 467
rect 1023 463 1057 467
rect 923 263 969 463
rect 1011 461 1069 463
rect 1017 458 1069 461
rect 994 453 1003 458
rect 1025 454 1069 458
rect 1082 454 1091 458
rect 983 442 1011 453
rect 1025 451 1063 454
rect 1023 442 1063 451
rect 994 275 1063 442
rect 1076 442 1091 454
rect 1103 454 1116 458
rect 994 266 1028 275
rect 994 263 1003 266
rect 1011 263 1026 266
rect 1040 263 1070 275
rect 935 259 948 263
rect 960 259 969 263
rect 982 259 1070 263
rect 939 254 1070 259
rect 1076 266 1095 442
rect 1076 254 1091 266
rect 994 250 1028 254
rect 967 225 1025 231
rect 1040 228 1070 254
rect 1082 250 1091 254
rect 1103 254 1128 454
rect 1137 254 1266 508
rect 1336 500 1394 506
rect 1336 466 1348 500
rect 1336 460 1394 466
rect 1103 250 1116 254
rect 880 177 909 225
rect 963 216 1029 225
rect 1137 216 1150 254
rect 967 210 979 216
rect 1154 210 1266 254
rect 963 191 1029 210
rect 967 185 1025 191
rect 1137 185 1266 210
rect 880 176 914 177
rect 880 142 1137 176
rect 846 108 1137 123
rect 1154 106 1266 185
rect 1336 172 1394 178
rect 1336 138 1348 172
rect 1336 132 1394 138
rect 1637 123 1646 603
rect 1671 517 1700 603
rect 1767 594 1925 603
rect 1671 225 1705 517
rect 1791 505 1804 535
rect 1820 526 1847 535
rect 1829 505 1842 526
rect 1945 508 2057 638
rect 1789 501 1816 505
rect 1817 501 1844 505
rect 1789 495 1879 501
rect 1813 492 1879 495
rect 1817 491 1844 492
rect 1817 486 1875 491
rect 1813 476 1844 485
rect 1831 467 1844 476
rect 1726 463 1739 467
rect 1751 463 1760 467
rect 1814 463 1848 467
rect 1714 263 1760 463
rect 1802 461 1860 463
rect 1808 458 1860 461
rect 1785 453 1794 458
rect 1816 454 1860 458
rect 1873 454 1882 458
rect 1774 442 1802 453
rect 1816 451 1854 454
rect 1814 442 1854 451
rect 1785 275 1854 442
rect 1867 442 1882 454
rect 1894 454 1907 458
rect 1785 266 1819 275
rect 1785 263 1794 266
rect 1802 263 1817 266
rect 1831 263 1861 275
rect 1726 259 1739 263
rect 1751 259 1760 263
rect 1773 259 1861 263
rect 1730 254 1861 259
rect 1867 266 1886 442
rect 1867 254 1882 266
rect 1785 250 1819 254
rect 1758 225 1816 231
rect 1831 228 1861 254
rect 1873 250 1882 254
rect 1894 254 1919 454
rect 1928 254 2057 508
rect 2127 500 2185 506
rect 2127 466 2139 500
rect 2127 460 2185 466
rect 1894 250 1907 254
rect 1671 177 1700 225
rect 1754 216 1820 225
rect 1928 216 1941 254
rect 1758 210 1770 216
rect 1945 210 2057 254
rect 1754 191 1820 210
rect 1758 185 1816 191
rect 1928 185 2057 210
rect 1671 176 1705 177
rect 1671 142 1928 176
rect 1637 108 1928 123
rect 1945 106 2057 185
rect 2127 172 2185 178
rect 2127 138 2139 172
rect 2127 132 2185 138
rect 363 89 433 106
rect 1154 89 1224 106
rect 1945 89 2015 106
rect 363 53 416 89
rect 1154 53 1207 89
rect 1945 53 1998 89
use inverter  x1
timestamp 1729033185
transform 1 0 -152 0 1 1
box 146 -1 937 1145
use inverter  x2
timestamp 1729033185
transform 1 0 639 0 1 1
box 146 -1 937 1145
use inverter  x3
timestamp 1729033185
transform 1 0 1430 0 1 1
box 146 -1 937 1145
<< end >>
