magic
tech sky130A
magscale 1 2
timestamp 1730269323
<< metal3 >>
rect -386 92012 386 92040
rect -386 91588 302 92012
rect 366 91588 386 92012
rect -386 91560 386 91588
rect -386 91292 386 91320
rect -386 90868 302 91292
rect 366 90868 386 91292
rect -386 90840 386 90868
rect -386 90572 386 90600
rect -386 90148 302 90572
rect 366 90148 386 90572
rect -386 90120 386 90148
rect -386 89852 386 89880
rect -386 89428 302 89852
rect 366 89428 386 89852
rect -386 89400 386 89428
rect -386 89132 386 89160
rect -386 88708 302 89132
rect 366 88708 386 89132
rect -386 88680 386 88708
rect -386 88412 386 88440
rect -386 87988 302 88412
rect 366 87988 386 88412
rect -386 87960 386 87988
rect -386 87692 386 87720
rect -386 87268 302 87692
rect 366 87268 386 87692
rect -386 87240 386 87268
rect -386 86972 386 87000
rect -386 86548 302 86972
rect 366 86548 386 86972
rect -386 86520 386 86548
rect -386 86252 386 86280
rect -386 85828 302 86252
rect 366 85828 386 86252
rect -386 85800 386 85828
rect -386 85532 386 85560
rect -386 85108 302 85532
rect 366 85108 386 85532
rect -386 85080 386 85108
rect -386 84812 386 84840
rect -386 84388 302 84812
rect 366 84388 386 84812
rect -386 84360 386 84388
rect -386 84092 386 84120
rect -386 83668 302 84092
rect 366 83668 386 84092
rect -386 83640 386 83668
rect -386 83372 386 83400
rect -386 82948 302 83372
rect 366 82948 386 83372
rect -386 82920 386 82948
rect -386 82652 386 82680
rect -386 82228 302 82652
rect 366 82228 386 82652
rect -386 82200 386 82228
rect -386 81932 386 81960
rect -386 81508 302 81932
rect 366 81508 386 81932
rect -386 81480 386 81508
rect -386 81212 386 81240
rect -386 80788 302 81212
rect 366 80788 386 81212
rect -386 80760 386 80788
rect -386 80492 386 80520
rect -386 80068 302 80492
rect 366 80068 386 80492
rect -386 80040 386 80068
rect -386 79772 386 79800
rect -386 79348 302 79772
rect 366 79348 386 79772
rect -386 79320 386 79348
rect -386 79052 386 79080
rect -386 78628 302 79052
rect 366 78628 386 79052
rect -386 78600 386 78628
rect -386 78332 386 78360
rect -386 77908 302 78332
rect 366 77908 386 78332
rect -386 77880 386 77908
rect -386 77612 386 77640
rect -386 77188 302 77612
rect 366 77188 386 77612
rect -386 77160 386 77188
rect -386 76892 386 76920
rect -386 76468 302 76892
rect 366 76468 386 76892
rect -386 76440 386 76468
rect -386 76172 386 76200
rect -386 75748 302 76172
rect 366 75748 386 76172
rect -386 75720 386 75748
rect -386 75452 386 75480
rect -386 75028 302 75452
rect 366 75028 386 75452
rect -386 75000 386 75028
rect -386 74732 386 74760
rect -386 74308 302 74732
rect 366 74308 386 74732
rect -386 74280 386 74308
rect -386 74012 386 74040
rect -386 73588 302 74012
rect 366 73588 386 74012
rect -386 73560 386 73588
rect -386 73292 386 73320
rect -386 72868 302 73292
rect 366 72868 386 73292
rect -386 72840 386 72868
rect -386 72572 386 72600
rect -386 72148 302 72572
rect 366 72148 386 72572
rect -386 72120 386 72148
rect -386 71852 386 71880
rect -386 71428 302 71852
rect 366 71428 386 71852
rect -386 71400 386 71428
rect -386 71132 386 71160
rect -386 70708 302 71132
rect 366 70708 386 71132
rect -386 70680 386 70708
rect -386 70412 386 70440
rect -386 69988 302 70412
rect 366 69988 386 70412
rect -386 69960 386 69988
rect -386 69692 386 69720
rect -386 69268 302 69692
rect 366 69268 386 69692
rect -386 69240 386 69268
rect -386 68972 386 69000
rect -386 68548 302 68972
rect 366 68548 386 68972
rect -386 68520 386 68548
rect -386 68252 386 68280
rect -386 67828 302 68252
rect 366 67828 386 68252
rect -386 67800 386 67828
rect -386 67532 386 67560
rect -386 67108 302 67532
rect 366 67108 386 67532
rect -386 67080 386 67108
rect -386 66812 386 66840
rect -386 66388 302 66812
rect 366 66388 386 66812
rect -386 66360 386 66388
rect -386 66092 386 66120
rect -386 65668 302 66092
rect 366 65668 386 66092
rect -386 65640 386 65668
rect -386 65372 386 65400
rect -386 64948 302 65372
rect 366 64948 386 65372
rect -386 64920 386 64948
rect -386 64652 386 64680
rect -386 64228 302 64652
rect 366 64228 386 64652
rect -386 64200 386 64228
rect -386 63932 386 63960
rect -386 63508 302 63932
rect 366 63508 386 63932
rect -386 63480 386 63508
rect -386 63212 386 63240
rect -386 62788 302 63212
rect 366 62788 386 63212
rect -386 62760 386 62788
rect -386 62492 386 62520
rect -386 62068 302 62492
rect 366 62068 386 62492
rect -386 62040 386 62068
rect -386 61772 386 61800
rect -386 61348 302 61772
rect 366 61348 386 61772
rect -386 61320 386 61348
rect -386 61052 386 61080
rect -386 60628 302 61052
rect 366 60628 386 61052
rect -386 60600 386 60628
rect -386 60332 386 60360
rect -386 59908 302 60332
rect 366 59908 386 60332
rect -386 59880 386 59908
rect -386 59612 386 59640
rect -386 59188 302 59612
rect 366 59188 386 59612
rect -386 59160 386 59188
rect -386 58892 386 58920
rect -386 58468 302 58892
rect 366 58468 386 58892
rect -386 58440 386 58468
rect -386 58172 386 58200
rect -386 57748 302 58172
rect 366 57748 386 58172
rect -386 57720 386 57748
rect -386 57452 386 57480
rect -386 57028 302 57452
rect 366 57028 386 57452
rect -386 57000 386 57028
rect -386 56732 386 56760
rect -386 56308 302 56732
rect 366 56308 386 56732
rect -386 56280 386 56308
rect -386 56012 386 56040
rect -386 55588 302 56012
rect 366 55588 386 56012
rect -386 55560 386 55588
rect -386 55292 386 55320
rect -386 54868 302 55292
rect 366 54868 386 55292
rect -386 54840 386 54868
rect -386 54572 386 54600
rect -386 54148 302 54572
rect 366 54148 386 54572
rect -386 54120 386 54148
rect -386 53852 386 53880
rect -386 53428 302 53852
rect 366 53428 386 53852
rect -386 53400 386 53428
rect -386 53132 386 53160
rect -386 52708 302 53132
rect 366 52708 386 53132
rect -386 52680 386 52708
rect -386 52412 386 52440
rect -386 51988 302 52412
rect 366 51988 386 52412
rect -386 51960 386 51988
rect -386 51692 386 51720
rect -386 51268 302 51692
rect 366 51268 386 51692
rect -386 51240 386 51268
rect -386 50972 386 51000
rect -386 50548 302 50972
rect 366 50548 386 50972
rect -386 50520 386 50548
rect -386 50252 386 50280
rect -386 49828 302 50252
rect 366 49828 386 50252
rect -386 49800 386 49828
rect -386 49532 386 49560
rect -386 49108 302 49532
rect 366 49108 386 49532
rect -386 49080 386 49108
rect -386 48812 386 48840
rect -386 48388 302 48812
rect 366 48388 386 48812
rect -386 48360 386 48388
rect -386 48092 386 48120
rect -386 47668 302 48092
rect 366 47668 386 48092
rect -386 47640 386 47668
rect -386 47372 386 47400
rect -386 46948 302 47372
rect 366 46948 386 47372
rect -386 46920 386 46948
rect -386 46652 386 46680
rect -386 46228 302 46652
rect 366 46228 386 46652
rect -386 46200 386 46228
rect -386 45932 386 45960
rect -386 45508 302 45932
rect 366 45508 386 45932
rect -386 45480 386 45508
rect -386 45212 386 45240
rect -386 44788 302 45212
rect 366 44788 386 45212
rect -386 44760 386 44788
rect -386 44492 386 44520
rect -386 44068 302 44492
rect 366 44068 386 44492
rect -386 44040 386 44068
rect -386 43772 386 43800
rect -386 43348 302 43772
rect 366 43348 386 43772
rect -386 43320 386 43348
rect -386 43052 386 43080
rect -386 42628 302 43052
rect 366 42628 386 43052
rect -386 42600 386 42628
rect -386 42332 386 42360
rect -386 41908 302 42332
rect 366 41908 386 42332
rect -386 41880 386 41908
rect -386 41612 386 41640
rect -386 41188 302 41612
rect 366 41188 386 41612
rect -386 41160 386 41188
rect -386 40892 386 40920
rect -386 40468 302 40892
rect 366 40468 386 40892
rect -386 40440 386 40468
rect -386 40172 386 40200
rect -386 39748 302 40172
rect 366 39748 386 40172
rect -386 39720 386 39748
rect -386 39452 386 39480
rect -386 39028 302 39452
rect 366 39028 386 39452
rect -386 39000 386 39028
rect -386 38732 386 38760
rect -386 38308 302 38732
rect 366 38308 386 38732
rect -386 38280 386 38308
rect -386 38012 386 38040
rect -386 37588 302 38012
rect 366 37588 386 38012
rect -386 37560 386 37588
rect -386 37292 386 37320
rect -386 36868 302 37292
rect 366 36868 386 37292
rect -386 36840 386 36868
rect -386 36572 386 36600
rect -386 36148 302 36572
rect 366 36148 386 36572
rect -386 36120 386 36148
rect -386 35852 386 35880
rect -386 35428 302 35852
rect 366 35428 386 35852
rect -386 35400 386 35428
rect -386 35132 386 35160
rect -386 34708 302 35132
rect 366 34708 386 35132
rect -386 34680 386 34708
rect -386 34412 386 34440
rect -386 33988 302 34412
rect 366 33988 386 34412
rect -386 33960 386 33988
rect -386 33692 386 33720
rect -386 33268 302 33692
rect 366 33268 386 33692
rect -386 33240 386 33268
rect -386 32972 386 33000
rect -386 32548 302 32972
rect 366 32548 386 32972
rect -386 32520 386 32548
rect -386 32252 386 32280
rect -386 31828 302 32252
rect 366 31828 386 32252
rect -386 31800 386 31828
rect -386 31532 386 31560
rect -386 31108 302 31532
rect 366 31108 386 31532
rect -386 31080 386 31108
rect -386 30812 386 30840
rect -386 30388 302 30812
rect 366 30388 386 30812
rect -386 30360 386 30388
rect -386 30092 386 30120
rect -386 29668 302 30092
rect 366 29668 386 30092
rect -386 29640 386 29668
rect -386 29372 386 29400
rect -386 28948 302 29372
rect 366 28948 386 29372
rect -386 28920 386 28948
rect -386 28652 386 28680
rect -386 28228 302 28652
rect 366 28228 386 28652
rect -386 28200 386 28228
rect -386 27932 386 27960
rect -386 27508 302 27932
rect 366 27508 386 27932
rect -386 27480 386 27508
rect -386 27212 386 27240
rect -386 26788 302 27212
rect 366 26788 386 27212
rect -386 26760 386 26788
rect -386 26492 386 26520
rect -386 26068 302 26492
rect 366 26068 386 26492
rect -386 26040 386 26068
rect -386 25772 386 25800
rect -386 25348 302 25772
rect 366 25348 386 25772
rect -386 25320 386 25348
rect -386 25052 386 25080
rect -386 24628 302 25052
rect 366 24628 386 25052
rect -386 24600 386 24628
rect -386 24332 386 24360
rect -386 23908 302 24332
rect 366 23908 386 24332
rect -386 23880 386 23908
rect -386 23612 386 23640
rect -386 23188 302 23612
rect 366 23188 386 23612
rect -386 23160 386 23188
rect -386 22892 386 22920
rect -386 22468 302 22892
rect 366 22468 386 22892
rect -386 22440 386 22468
rect -386 22172 386 22200
rect -386 21748 302 22172
rect 366 21748 386 22172
rect -386 21720 386 21748
rect -386 21452 386 21480
rect -386 21028 302 21452
rect 366 21028 386 21452
rect -386 21000 386 21028
rect -386 20732 386 20760
rect -386 20308 302 20732
rect 366 20308 386 20732
rect -386 20280 386 20308
rect -386 20012 386 20040
rect -386 19588 302 20012
rect 366 19588 386 20012
rect -386 19560 386 19588
rect -386 19292 386 19320
rect -386 18868 302 19292
rect 366 18868 386 19292
rect -386 18840 386 18868
rect -386 18572 386 18600
rect -386 18148 302 18572
rect 366 18148 386 18572
rect -386 18120 386 18148
rect -386 17852 386 17880
rect -386 17428 302 17852
rect 366 17428 386 17852
rect -386 17400 386 17428
rect -386 17132 386 17160
rect -386 16708 302 17132
rect 366 16708 386 17132
rect -386 16680 386 16708
rect -386 16412 386 16440
rect -386 15988 302 16412
rect 366 15988 386 16412
rect -386 15960 386 15988
rect -386 15692 386 15720
rect -386 15268 302 15692
rect 366 15268 386 15692
rect -386 15240 386 15268
rect -386 14972 386 15000
rect -386 14548 302 14972
rect 366 14548 386 14972
rect -386 14520 386 14548
rect -386 14252 386 14280
rect -386 13828 302 14252
rect 366 13828 386 14252
rect -386 13800 386 13828
rect -386 13532 386 13560
rect -386 13108 302 13532
rect 366 13108 386 13532
rect -386 13080 386 13108
rect -386 12812 386 12840
rect -386 12388 302 12812
rect 366 12388 386 12812
rect -386 12360 386 12388
rect -386 12092 386 12120
rect -386 11668 302 12092
rect 366 11668 386 12092
rect -386 11640 386 11668
rect -386 11372 386 11400
rect -386 10948 302 11372
rect 366 10948 386 11372
rect -386 10920 386 10948
rect -386 10652 386 10680
rect -386 10228 302 10652
rect 366 10228 386 10652
rect -386 10200 386 10228
rect -386 9932 386 9960
rect -386 9508 302 9932
rect 366 9508 386 9932
rect -386 9480 386 9508
rect -386 9212 386 9240
rect -386 8788 302 9212
rect 366 8788 386 9212
rect -386 8760 386 8788
rect -386 8492 386 8520
rect -386 8068 302 8492
rect 366 8068 386 8492
rect -386 8040 386 8068
rect -386 7772 386 7800
rect -386 7348 302 7772
rect 366 7348 386 7772
rect -386 7320 386 7348
rect -386 7052 386 7080
rect -386 6628 302 7052
rect 366 6628 386 7052
rect -386 6600 386 6628
rect -386 6332 386 6360
rect -386 5908 302 6332
rect 366 5908 386 6332
rect -386 5880 386 5908
rect -386 5612 386 5640
rect -386 5188 302 5612
rect 366 5188 386 5612
rect -386 5160 386 5188
rect -386 4892 386 4920
rect -386 4468 302 4892
rect 366 4468 386 4892
rect -386 4440 386 4468
rect -386 4172 386 4200
rect -386 3748 302 4172
rect 366 3748 386 4172
rect -386 3720 386 3748
rect -386 3452 386 3480
rect -386 3028 302 3452
rect 366 3028 386 3452
rect -386 3000 386 3028
rect -386 2732 386 2760
rect -386 2308 302 2732
rect 366 2308 386 2732
rect -386 2280 386 2308
rect -386 2012 386 2040
rect -386 1588 302 2012
rect 366 1588 386 2012
rect -386 1560 386 1588
rect -386 1292 386 1320
rect -386 868 302 1292
rect 366 868 386 1292
rect -386 840 386 868
rect -386 572 386 600
rect -386 148 302 572
rect 366 148 386 572
rect -386 120 386 148
rect -386 -148 386 -120
rect -386 -572 302 -148
rect 366 -572 386 -148
rect -386 -600 386 -572
rect -386 -868 386 -840
rect -386 -1292 302 -868
rect 366 -1292 386 -868
rect -386 -1320 386 -1292
rect -386 -1588 386 -1560
rect -386 -2012 302 -1588
rect 366 -2012 386 -1588
rect -386 -2040 386 -2012
rect -386 -2308 386 -2280
rect -386 -2732 302 -2308
rect 366 -2732 386 -2308
rect -386 -2760 386 -2732
rect -386 -3028 386 -3000
rect -386 -3452 302 -3028
rect 366 -3452 386 -3028
rect -386 -3480 386 -3452
rect -386 -3748 386 -3720
rect -386 -4172 302 -3748
rect 366 -4172 386 -3748
rect -386 -4200 386 -4172
rect -386 -4468 386 -4440
rect -386 -4892 302 -4468
rect 366 -4892 386 -4468
rect -386 -4920 386 -4892
rect -386 -5188 386 -5160
rect -386 -5612 302 -5188
rect 366 -5612 386 -5188
rect -386 -5640 386 -5612
rect -386 -5908 386 -5880
rect -386 -6332 302 -5908
rect 366 -6332 386 -5908
rect -386 -6360 386 -6332
rect -386 -6628 386 -6600
rect -386 -7052 302 -6628
rect 366 -7052 386 -6628
rect -386 -7080 386 -7052
rect -386 -7348 386 -7320
rect -386 -7772 302 -7348
rect 366 -7772 386 -7348
rect -386 -7800 386 -7772
rect -386 -8068 386 -8040
rect -386 -8492 302 -8068
rect 366 -8492 386 -8068
rect -386 -8520 386 -8492
rect -386 -8788 386 -8760
rect -386 -9212 302 -8788
rect 366 -9212 386 -8788
rect -386 -9240 386 -9212
rect -386 -9508 386 -9480
rect -386 -9932 302 -9508
rect 366 -9932 386 -9508
rect -386 -9960 386 -9932
rect -386 -10228 386 -10200
rect -386 -10652 302 -10228
rect 366 -10652 386 -10228
rect -386 -10680 386 -10652
rect -386 -10948 386 -10920
rect -386 -11372 302 -10948
rect 366 -11372 386 -10948
rect -386 -11400 386 -11372
rect -386 -11668 386 -11640
rect -386 -12092 302 -11668
rect 366 -12092 386 -11668
rect -386 -12120 386 -12092
rect -386 -12388 386 -12360
rect -386 -12812 302 -12388
rect 366 -12812 386 -12388
rect -386 -12840 386 -12812
rect -386 -13108 386 -13080
rect -386 -13532 302 -13108
rect 366 -13532 386 -13108
rect -386 -13560 386 -13532
rect -386 -13828 386 -13800
rect -386 -14252 302 -13828
rect 366 -14252 386 -13828
rect -386 -14280 386 -14252
rect -386 -14548 386 -14520
rect -386 -14972 302 -14548
rect 366 -14972 386 -14548
rect -386 -15000 386 -14972
rect -386 -15268 386 -15240
rect -386 -15692 302 -15268
rect 366 -15692 386 -15268
rect -386 -15720 386 -15692
rect -386 -15988 386 -15960
rect -386 -16412 302 -15988
rect 366 -16412 386 -15988
rect -386 -16440 386 -16412
rect -386 -16708 386 -16680
rect -386 -17132 302 -16708
rect 366 -17132 386 -16708
rect -386 -17160 386 -17132
rect -386 -17428 386 -17400
rect -386 -17852 302 -17428
rect 366 -17852 386 -17428
rect -386 -17880 386 -17852
rect -386 -18148 386 -18120
rect -386 -18572 302 -18148
rect 366 -18572 386 -18148
rect -386 -18600 386 -18572
rect -386 -18868 386 -18840
rect -386 -19292 302 -18868
rect 366 -19292 386 -18868
rect -386 -19320 386 -19292
rect -386 -19588 386 -19560
rect -386 -20012 302 -19588
rect 366 -20012 386 -19588
rect -386 -20040 386 -20012
rect -386 -20308 386 -20280
rect -386 -20732 302 -20308
rect 366 -20732 386 -20308
rect -386 -20760 386 -20732
rect -386 -21028 386 -21000
rect -386 -21452 302 -21028
rect 366 -21452 386 -21028
rect -386 -21480 386 -21452
rect -386 -21748 386 -21720
rect -386 -22172 302 -21748
rect 366 -22172 386 -21748
rect -386 -22200 386 -22172
rect -386 -22468 386 -22440
rect -386 -22892 302 -22468
rect 366 -22892 386 -22468
rect -386 -22920 386 -22892
rect -386 -23188 386 -23160
rect -386 -23612 302 -23188
rect 366 -23612 386 -23188
rect -386 -23640 386 -23612
rect -386 -23908 386 -23880
rect -386 -24332 302 -23908
rect 366 -24332 386 -23908
rect -386 -24360 386 -24332
rect -386 -24628 386 -24600
rect -386 -25052 302 -24628
rect 366 -25052 386 -24628
rect -386 -25080 386 -25052
rect -386 -25348 386 -25320
rect -386 -25772 302 -25348
rect 366 -25772 386 -25348
rect -386 -25800 386 -25772
rect -386 -26068 386 -26040
rect -386 -26492 302 -26068
rect 366 -26492 386 -26068
rect -386 -26520 386 -26492
rect -386 -26788 386 -26760
rect -386 -27212 302 -26788
rect 366 -27212 386 -26788
rect -386 -27240 386 -27212
rect -386 -27508 386 -27480
rect -386 -27932 302 -27508
rect 366 -27932 386 -27508
rect -386 -27960 386 -27932
rect -386 -28228 386 -28200
rect -386 -28652 302 -28228
rect 366 -28652 386 -28228
rect -386 -28680 386 -28652
rect -386 -28948 386 -28920
rect -386 -29372 302 -28948
rect 366 -29372 386 -28948
rect -386 -29400 386 -29372
rect -386 -29668 386 -29640
rect -386 -30092 302 -29668
rect 366 -30092 386 -29668
rect -386 -30120 386 -30092
rect -386 -30388 386 -30360
rect -386 -30812 302 -30388
rect 366 -30812 386 -30388
rect -386 -30840 386 -30812
rect -386 -31108 386 -31080
rect -386 -31532 302 -31108
rect 366 -31532 386 -31108
rect -386 -31560 386 -31532
rect -386 -31828 386 -31800
rect -386 -32252 302 -31828
rect 366 -32252 386 -31828
rect -386 -32280 386 -32252
rect -386 -32548 386 -32520
rect -386 -32972 302 -32548
rect 366 -32972 386 -32548
rect -386 -33000 386 -32972
rect -386 -33268 386 -33240
rect -386 -33692 302 -33268
rect 366 -33692 386 -33268
rect -386 -33720 386 -33692
rect -386 -33988 386 -33960
rect -386 -34412 302 -33988
rect 366 -34412 386 -33988
rect -386 -34440 386 -34412
rect -386 -34708 386 -34680
rect -386 -35132 302 -34708
rect 366 -35132 386 -34708
rect -386 -35160 386 -35132
rect -386 -35428 386 -35400
rect -386 -35852 302 -35428
rect 366 -35852 386 -35428
rect -386 -35880 386 -35852
rect -386 -36148 386 -36120
rect -386 -36572 302 -36148
rect 366 -36572 386 -36148
rect -386 -36600 386 -36572
rect -386 -36868 386 -36840
rect -386 -37292 302 -36868
rect 366 -37292 386 -36868
rect -386 -37320 386 -37292
rect -386 -37588 386 -37560
rect -386 -38012 302 -37588
rect 366 -38012 386 -37588
rect -386 -38040 386 -38012
rect -386 -38308 386 -38280
rect -386 -38732 302 -38308
rect 366 -38732 386 -38308
rect -386 -38760 386 -38732
rect -386 -39028 386 -39000
rect -386 -39452 302 -39028
rect 366 -39452 386 -39028
rect -386 -39480 386 -39452
rect -386 -39748 386 -39720
rect -386 -40172 302 -39748
rect 366 -40172 386 -39748
rect -386 -40200 386 -40172
rect -386 -40468 386 -40440
rect -386 -40892 302 -40468
rect 366 -40892 386 -40468
rect -386 -40920 386 -40892
rect -386 -41188 386 -41160
rect -386 -41612 302 -41188
rect 366 -41612 386 -41188
rect -386 -41640 386 -41612
rect -386 -41908 386 -41880
rect -386 -42332 302 -41908
rect 366 -42332 386 -41908
rect -386 -42360 386 -42332
rect -386 -42628 386 -42600
rect -386 -43052 302 -42628
rect 366 -43052 386 -42628
rect -386 -43080 386 -43052
rect -386 -43348 386 -43320
rect -386 -43772 302 -43348
rect 366 -43772 386 -43348
rect -386 -43800 386 -43772
rect -386 -44068 386 -44040
rect -386 -44492 302 -44068
rect 366 -44492 386 -44068
rect -386 -44520 386 -44492
rect -386 -44788 386 -44760
rect -386 -45212 302 -44788
rect 366 -45212 386 -44788
rect -386 -45240 386 -45212
rect -386 -45508 386 -45480
rect -386 -45932 302 -45508
rect 366 -45932 386 -45508
rect -386 -45960 386 -45932
rect -386 -46228 386 -46200
rect -386 -46652 302 -46228
rect 366 -46652 386 -46228
rect -386 -46680 386 -46652
rect -386 -46948 386 -46920
rect -386 -47372 302 -46948
rect 366 -47372 386 -46948
rect -386 -47400 386 -47372
rect -386 -47668 386 -47640
rect -386 -48092 302 -47668
rect 366 -48092 386 -47668
rect -386 -48120 386 -48092
rect -386 -48388 386 -48360
rect -386 -48812 302 -48388
rect 366 -48812 386 -48388
rect -386 -48840 386 -48812
rect -386 -49108 386 -49080
rect -386 -49532 302 -49108
rect 366 -49532 386 -49108
rect -386 -49560 386 -49532
rect -386 -49828 386 -49800
rect -386 -50252 302 -49828
rect 366 -50252 386 -49828
rect -386 -50280 386 -50252
rect -386 -50548 386 -50520
rect -386 -50972 302 -50548
rect 366 -50972 386 -50548
rect -386 -51000 386 -50972
rect -386 -51268 386 -51240
rect -386 -51692 302 -51268
rect 366 -51692 386 -51268
rect -386 -51720 386 -51692
rect -386 -51988 386 -51960
rect -386 -52412 302 -51988
rect 366 -52412 386 -51988
rect -386 -52440 386 -52412
rect -386 -52708 386 -52680
rect -386 -53132 302 -52708
rect 366 -53132 386 -52708
rect -386 -53160 386 -53132
rect -386 -53428 386 -53400
rect -386 -53852 302 -53428
rect 366 -53852 386 -53428
rect -386 -53880 386 -53852
rect -386 -54148 386 -54120
rect -386 -54572 302 -54148
rect 366 -54572 386 -54148
rect -386 -54600 386 -54572
rect -386 -54868 386 -54840
rect -386 -55292 302 -54868
rect 366 -55292 386 -54868
rect -386 -55320 386 -55292
rect -386 -55588 386 -55560
rect -386 -56012 302 -55588
rect 366 -56012 386 -55588
rect -386 -56040 386 -56012
rect -386 -56308 386 -56280
rect -386 -56732 302 -56308
rect 366 -56732 386 -56308
rect -386 -56760 386 -56732
rect -386 -57028 386 -57000
rect -386 -57452 302 -57028
rect 366 -57452 386 -57028
rect -386 -57480 386 -57452
rect -386 -57748 386 -57720
rect -386 -58172 302 -57748
rect 366 -58172 386 -57748
rect -386 -58200 386 -58172
rect -386 -58468 386 -58440
rect -386 -58892 302 -58468
rect 366 -58892 386 -58468
rect -386 -58920 386 -58892
rect -386 -59188 386 -59160
rect -386 -59612 302 -59188
rect 366 -59612 386 -59188
rect -386 -59640 386 -59612
rect -386 -59908 386 -59880
rect -386 -60332 302 -59908
rect 366 -60332 386 -59908
rect -386 -60360 386 -60332
rect -386 -60628 386 -60600
rect -386 -61052 302 -60628
rect 366 -61052 386 -60628
rect -386 -61080 386 -61052
rect -386 -61348 386 -61320
rect -386 -61772 302 -61348
rect 366 -61772 386 -61348
rect -386 -61800 386 -61772
rect -386 -62068 386 -62040
rect -386 -62492 302 -62068
rect 366 -62492 386 -62068
rect -386 -62520 386 -62492
rect -386 -62788 386 -62760
rect -386 -63212 302 -62788
rect 366 -63212 386 -62788
rect -386 -63240 386 -63212
rect -386 -63508 386 -63480
rect -386 -63932 302 -63508
rect 366 -63932 386 -63508
rect -386 -63960 386 -63932
rect -386 -64228 386 -64200
rect -386 -64652 302 -64228
rect 366 -64652 386 -64228
rect -386 -64680 386 -64652
rect -386 -64948 386 -64920
rect -386 -65372 302 -64948
rect 366 -65372 386 -64948
rect -386 -65400 386 -65372
rect -386 -65668 386 -65640
rect -386 -66092 302 -65668
rect 366 -66092 386 -65668
rect -386 -66120 386 -66092
rect -386 -66388 386 -66360
rect -386 -66812 302 -66388
rect 366 -66812 386 -66388
rect -386 -66840 386 -66812
rect -386 -67108 386 -67080
rect -386 -67532 302 -67108
rect 366 -67532 386 -67108
rect -386 -67560 386 -67532
rect -386 -67828 386 -67800
rect -386 -68252 302 -67828
rect 366 -68252 386 -67828
rect -386 -68280 386 -68252
rect -386 -68548 386 -68520
rect -386 -68972 302 -68548
rect 366 -68972 386 -68548
rect -386 -69000 386 -68972
rect -386 -69268 386 -69240
rect -386 -69692 302 -69268
rect 366 -69692 386 -69268
rect -386 -69720 386 -69692
rect -386 -69988 386 -69960
rect -386 -70412 302 -69988
rect 366 -70412 386 -69988
rect -386 -70440 386 -70412
rect -386 -70708 386 -70680
rect -386 -71132 302 -70708
rect 366 -71132 386 -70708
rect -386 -71160 386 -71132
rect -386 -71428 386 -71400
rect -386 -71852 302 -71428
rect 366 -71852 386 -71428
rect -386 -71880 386 -71852
rect -386 -72148 386 -72120
rect -386 -72572 302 -72148
rect 366 -72572 386 -72148
rect -386 -72600 386 -72572
rect -386 -72868 386 -72840
rect -386 -73292 302 -72868
rect 366 -73292 386 -72868
rect -386 -73320 386 -73292
rect -386 -73588 386 -73560
rect -386 -74012 302 -73588
rect 366 -74012 386 -73588
rect -386 -74040 386 -74012
rect -386 -74308 386 -74280
rect -386 -74732 302 -74308
rect 366 -74732 386 -74308
rect -386 -74760 386 -74732
rect -386 -75028 386 -75000
rect -386 -75452 302 -75028
rect 366 -75452 386 -75028
rect -386 -75480 386 -75452
rect -386 -75748 386 -75720
rect -386 -76172 302 -75748
rect 366 -76172 386 -75748
rect -386 -76200 386 -76172
rect -386 -76468 386 -76440
rect -386 -76892 302 -76468
rect 366 -76892 386 -76468
rect -386 -76920 386 -76892
rect -386 -77188 386 -77160
rect -386 -77612 302 -77188
rect 366 -77612 386 -77188
rect -386 -77640 386 -77612
rect -386 -77908 386 -77880
rect -386 -78332 302 -77908
rect 366 -78332 386 -77908
rect -386 -78360 386 -78332
rect -386 -78628 386 -78600
rect -386 -79052 302 -78628
rect 366 -79052 386 -78628
rect -386 -79080 386 -79052
rect -386 -79348 386 -79320
rect -386 -79772 302 -79348
rect 366 -79772 386 -79348
rect -386 -79800 386 -79772
rect -386 -80068 386 -80040
rect -386 -80492 302 -80068
rect 366 -80492 386 -80068
rect -386 -80520 386 -80492
rect -386 -80788 386 -80760
rect -386 -81212 302 -80788
rect 366 -81212 386 -80788
rect -386 -81240 386 -81212
rect -386 -81508 386 -81480
rect -386 -81932 302 -81508
rect 366 -81932 386 -81508
rect -386 -81960 386 -81932
rect -386 -82228 386 -82200
rect -386 -82652 302 -82228
rect 366 -82652 386 -82228
rect -386 -82680 386 -82652
rect -386 -82948 386 -82920
rect -386 -83372 302 -82948
rect 366 -83372 386 -82948
rect -386 -83400 386 -83372
rect -386 -83668 386 -83640
rect -386 -84092 302 -83668
rect 366 -84092 386 -83668
rect -386 -84120 386 -84092
rect -386 -84388 386 -84360
rect -386 -84812 302 -84388
rect 366 -84812 386 -84388
rect -386 -84840 386 -84812
rect -386 -85108 386 -85080
rect -386 -85532 302 -85108
rect 366 -85532 386 -85108
rect -386 -85560 386 -85532
rect -386 -85828 386 -85800
rect -386 -86252 302 -85828
rect 366 -86252 386 -85828
rect -386 -86280 386 -86252
rect -386 -86548 386 -86520
rect -386 -86972 302 -86548
rect 366 -86972 386 -86548
rect -386 -87000 386 -86972
rect -386 -87268 386 -87240
rect -386 -87692 302 -87268
rect 366 -87692 386 -87268
rect -386 -87720 386 -87692
rect -386 -87988 386 -87960
rect -386 -88412 302 -87988
rect 366 -88412 386 -87988
rect -386 -88440 386 -88412
rect -386 -88708 386 -88680
rect -386 -89132 302 -88708
rect 366 -89132 386 -88708
rect -386 -89160 386 -89132
rect -386 -89428 386 -89400
rect -386 -89852 302 -89428
rect 366 -89852 386 -89428
rect -386 -89880 386 -89852
rect -386 -90148 386 -90120
rect -386 -90572 302 -90148
rect 366 -90572 386 -90148
rect -386 -90600 386 -90572
rect -386 -90868 386 -90840
rect -386 -91292 302 -90868
rect 366 -91292 386 -90868
rect -386 -91320 386 -91292
rect -386 -91588 386 -91560
rect -386 -92012 302 -91588
rect 366 -92012 386 -91588
rect -386 -92040 386 -92012
<< via3 >>
rect 302 91588 366 92012
rect 302 90868 366 91292
rect 302 90148 366 90572
rect 302 89428 366 89852
rect 302 88708 366 89132
rect 302 87988 366 88412
rect 302 87268 366 87692
rect 302 86548 366 86972
rect 302 85828 366 86252
rect 302 85108 366 85532
rect 302 84388 366 84812
rect 302 83668 366 84092
rect 302 82948 366 83372
rect 302 82228 366 82652
rect 302 81508 366 81932
rect 302 80788 366 81212
rect 302 80068 366 80492
rect 302 79348 366 79772
rect 302 78628 366 79052
rect 302 77908 366 78332
rect 302 77188 366 77612
rect 302 76468 366 76892
rect 302 75748 366 76172
rect 302 75028 366 75452
rect 302 74308 366 74732
rect 302 73588 366 74012
rect 302 72868 366 73292
rect 302 72148 366 72572
rect 302 71428 366 71852
rect 302 70708 366 71132
rect 302 69988 366 70412
rect 302 69268 366 69692
rect 302 68548 366 68972
rect 302 67828 366 68252
rect 302 67108 366 67532
rect 302 66388 366 66812
rect 302 65668 366 66092
rect 302 64948 366 65372
rect 302 64228 366 64652
rect 302 63508 366 63932
rect 302 62788 366 63212
rect 302 62068 366 62492
rect 302 61348 366 61772
rect 302 60628 366 61052
rect 302 59908 366 60332
rect 302 59188 366 59612
rect 302 58468 366 58892
rect 302 57748 366 58172
rect 302 57028 366 57452
rect 302 56308 366 56732
rect 302 55588 366 56012
rect 302 54868 366 55292
rect 302 54148 366 54572
rect 302 53428 366 53852
rect 302 52708 366 53132
rect 302 51988 366 52412
rect 302 51268 366 51692
rect 302 50548 366 50972
rect 302 49828 366 50252
rect 302 49108 366 49532
rect 302 48388 366 48812
rect 302 47668 366 48092
rect 302 46948 366 47372
rect 302 46228 366 46652
rect 302 45508 366 45932
rect 302 44788 366 45212
rect 302 44068 366 44492
rect 302 43348 366 43772
rect 302 42628 366 43052
rect 302 41908 366 42332
rect 302 41188 366 41612
rect 302 40468 366 40892
rect 302 39748 366 40172
rect 302 39028 366 39452
rect 302 38308 366 38732
rect 302 37588 366 38012
rect 302 36868 366 37292
rect 302 36148 366 36572
rect 302 35428 366 35852
rect 302 34708 366 35132
rect 302 33988 366 34412
rect 302 33268 366 33692
rect 302 32548 366 32972
rect 302 31828 366 32252
rect 302 31108 366 31532
rect 302 30388 366 30812
rect 302 29668 366 30092
rect 302 28948 366 29372
rect 302 28228 366 28652
rect 302 27508 366 27932
rect 302 26788 366 27212
rect 302 26068 366 26492
rect 302 25348 366 25772
rect 302 24628 366 25052
rect 302 23908 366 24332
rect 302 23188 366 23612
rect 302 22468 366 22892
rect 302 21748 366 22172
rect 302 21028 366 21452
rect 302 20308 366 20732
rect 302 19588 366 20012
rect 302 18868 366 19292
rect 302 18148 366 18572
rect 302 17428 366 17852
rect 302 16708 366 17132
rect 302 15988 366 16412
rect 302 15268 366 15692
rect 302 14548 366 14972
rect 302 13828 366 14252
rect 302 13108 366 13532
rect 302 12388 366 12812
rect 302 11668 366 12092
rect 302 10948 366 11372
rect 302 10228 366 10652
rect 302 9508 366 9932
rect 302 8788 366 9212
rect 302 8068 366 8492
rect 302 7348 366 7772
rect 302 6628 366 7052
rect 302 5908 366 6332
rect 302 5188 366 5612
rect 302 4468 366 4892
rect 302 3748 366 4172
rect 302 3028 366 3452
rect 302 2308 366 2732
rect 302 1588 366 2012
rect 302 868 366 1292
rect 302 148 366 572
rect 302 -572 366 -148
rect 302 -1292 366 -868
rect 302 -2012 366 -1588
rect 302 -2732 366 -2308
rect 302 -3452 366 -3028
rect 302 -4172 366 -3748
rect 302 -4892 366 -4468
rect 302 -5612 366 -5188
rect 302 -6332 366 -5908
rect 302 -7052 366 -6628
rect 302 -7772 366 -7348
rect 302 -8492 366 -8068
rect 302 -9212 366 -8788
rect 302 -9932 366 -9508
rect 302 -10652 366 -10228
rect 302 -11372 366 -10948
rect 302 -12092 366 -11668
rect 302 -12812 366 -12388
rect 302 -13532 366 -13108
rect 302 -14252 366 -13828
rect 302 -14972 366 -14548
rect 302 -15692 366 -15268
rect 302 -16412 366 -15988
rect 302 -17132 366 -16708
rect 302 -17852 366 -17428
rect 302 -18572 366 -18148
rect 302 -19292 366 -18868
rect 302 -20012 366 -19588
rect 302 -20732 366 -20308
rect 302 -21452 366 -21028
rect 302 -22172 366 -21748
rect 302 -22892 366 -22468
rect 302 -23612 366 -23188
rect 302 -24332 366 -23908
rect 302 -25052 366 -24628
rect 302 -25772 366 -25348
rect 302 -26492 366 -26068
rect 302 -27212 366 -26788
rect 302 -27932 366 -27508
rect 302 -28652 366 -28228
rect 302 -29372 366 -28948
rect 302 -30092 366 -29668
rect 302 -30812 366 -30388
rect 302 -31532 366 -31108
rect 302 -32252 366 -31828
rect 302 -32972 366 -32548
rect 302 -33692 366 -33268
rect 302 -34412 366 -33988
rect 302 -35132 366 -34708
rect 302 -35852 366 -35428
rect 302 -36572 366 -36148
rect 302 -37292 366 -36868
rect 302 -38012 366 -37588
rect 302 -38732 366 -38308
rect 302 -39452 366 -39028
rect 302 -40172 366 -39748
rect 302 -40892 366 -40468
rect 302 -41612 366 -41188
rect 302 -42332 366 -41908
rect 302 -43052 366 -42628
rect 302 -43772 366 -43348
rect 302 -44492 366 -44068
rect 302 -45212 366 -44788
rect 302 -45932 366 -45508
rect 302 -46652 366 -46228
rect 302 -47372 366 -46948
rect 302 -48092 366 -47668
rect 302 -48812 366 -48388
rect 302 -49532 366 -49108
rect 302 -50252 366 -49828
rect 302 -50972 366 -50548
rect 302 -51692 366 -51268
rect 302 -52412 366 -51988
rect 302 -53132 366 -52708
rect 302 -53852 366 -53428
rect 302 -54572 366 -54148
rect 302 -55292 366 -54868
rect 302 -56012 366 -55588
rect 302 -56732 366 -56308
rect 302 -57452 366 -57028
rect 302 -58172 366 -57748
rect 302 -58892 366 -58468
rect 302 -59612 366 -59188
rect 302 -60332 366 -59908
rect 302 -61052 366 -60628
rect 302 -61772 366 -61348
rect 302 -62492 366 -62068
rect 302 -63212 366 -62788
rect 302 -63932 366 -63508
rect 302 -64652 366 -64228
rect 302 -65372 366 -64948
rect 302 -66092 366 -65668
rect 302 -66812 366 -66388
rect 302 -67532 366 -67108
rect 302 -68252 366 -67828
rect 302 -68972 366 -68548
rect 302 -69692 366 -69268
rect 302 -70412 366 -69988
rect 302 -71132 366 -70708
rect 302 -71852 366 -71428
rect 302 -72572 366 -72148
rect 302 -73292 366 -72868
rect 302 -74012 366 -73588
rect 302 -74732 366 -74308
rect 302 -75452 366 -75028
rect 302 -76172 366 -75748
rect 302 -76892 366 -76468
rect 302 -77612 366 -77188
rect 302 -78332 366 -77908
rect 302 -79052 366 -78628
rect 302 -79772 366 -79348
rect 302 -80492 366 -80068
rect 302 -81212 366 -80788
rect 302 -81932 366 -81508
rect 302 -82652 366 -82228
rect 302 -83372 366 -82948
rect 302 -84092 366 -83668
rect 302 -84812 366 -84388
rect 302 -85532 366 -85108
rect 302 -86252 366 -85828
rect 302 -86972 366 -86548
rect 302 -87692 366 -87268
rect 302 -88412 366 -87988
rect 302 -89132 366 -88708
rect 302 -89852 366 -89428
rect 302 -90572 366 -90148
rect 302 -91292 366 -90868
rect 302 -92012 366 -91588
<< mimcap >>
rect -346 91960 54 92000
rect -346 91640 -306 91960
rect 14 91640 54 91960
rect -346 91600 54 91640
rect -346 91240 54 91280
rect -346 90920 -306 91240
rect 14 90920 54 91240
rect -346 90880 54 90920
rect -346 90520 54 90560
rect -346 90200 -306 90520
rect 14 90200 54 90520
rect -346 90160 54 90200
rect -346 89800 54 89840
rect -346 89480 -306 89800
rect 14 89480 54 89800
rect -346 89440 54 89480
rect -346 89080 54 89120
rect -346 88760 -306 89080
rect 14 88760 54 89080
rect -346 88720 54 88760
rect -346 88360 54 88400
rect -346 88040 -306 88360
rect 14 88040 54 88360
rect -346 88000 54 88040
rect -346 87640 54 87680
rect -346 87320 -306 87640
rect 14 87320 54 87640
rect -346 87280 54 87320
rect -346 86920 54 86960
rect -346 86600 -306 86920
rect 14 86600 54 86920
rect -346 86560 54 86600
rect -346 86200 54 86240
rect -346 85880 -306 86200
rect 14 85880 54 86200
rect -346 85840 54 85880
rect -346 85480 54 85520
rect -346 85160 -306 85480
rect 14 85160 54 85480
rect -346 85120 54 85160
rect -346 84760 54 84800
rect -346 84440 -306 84760
rect 14 84440 54 84760
rect -346 84400 54 84440
rect -346 84040 54 84080
rect -346 83720 -306 84040
rect 14 83720 54 84040
rect -346 83680 54 83720
rect -346 83320 54 83360
rect -346 83000 -306 83320
rect 14 83000 54 83320
rect -346 82960 54 83000
rect -346 82600 54 82640
rect -346 82280 -306 82600
rect 14 82280 54 82600
rect -346 82240 54 82280
rect -346 81880 54 81920
rect -346 81560 -306 81880
rect 14 81560 54 81880
rect -346 81520 54 81560
rect -346 81160 54 81200
rect -346 80840 -306 81160
rect 14 80840 54 81160
rect -346 80800 54 80840
rect -346 80440 54 80480
rect -346 80120 -306 80440
rect 14 80120 54 80440
rect -346 80080 54 80120
rect -346 79720 54 79760
rect -346 79400 -306 79720
rect 14 79400 54 79720
rect -346 79360 54 79400
rect -346 79000 54 79040
rect -346 78680 -306 79000
rect 14 78680 54 79000
rect -346 78640 54 78680
rect -346 78280 54 78320
rect -346 77960 -306 78280
rect 14 77960 54 78280
rect -346 77920 54 77960
rect -346 77560 54 77600
rect -346 77240 -306 77560
rect 14 77240 54 77560
rect -346 77200 54 77240
rect -346 76840 54 76880
rect -346 76520 -306 76840
rect 14 76520 54 76840
rect -346 76480 54 76520
rect -346 76120 54 76160
rect -346 75800 -306 76120
rect 14 75800 54 76120
rect -346 75760 54 75800
rect -346 75400 54 75440
rect -346 75080 -306 75400
rect 14 75080 54 75400
rect -346 75040 54 75080
rect -346 74680 54 74720
rect -346 74360 -306 74680
rect 14 74360 54 74680
rect -346 74320 54 74360
rect -346 73960 54 74000
rect -346 73640 -306 73960
rect 14 73640 54 73960
rect -346 73600 54 73640
rect -346 73240 54 73280
rect -346 72920 -306 73240
rect 14 72920 54 73240
rect -346 72880 54 72920
rect -346 72520 54 72560
rect -346 72200 -306 72520
rect 14 72200 54 72520
rect -346 72160 54 72200
rect -346 71800 54 71840
rect -346 71480 -306 71800
rect 14 71480 54 71800
rect -346 71440 54 71480
rect -346 71080 54 71120
rect -346 70760 -306 71080
rect 14 70760 54 71080
rect -346 70720 54 70760
rect -346 70360 54 70400
rect -346 70040 -306 70360
rect 14 70040 54 70360
rect -346 70000 54 70040
rect -346 69640 54 69680
rect -346 69320 -306 69640
rect 14 69320 54 69640
rect -346 69280 54 69320
rect -346 68920 54 68960
rect -346 68600 -306 68920
rect 14 68600 54 68920
rect -346 68560 54 68600
rect -346 68200 54 68240
rect -346 67880 -306 68200
rect 14 67880 54 68200
rect -346 67840 54 67880
rect -346 67480 54 67520
rect -346 67160 -306 67480
rect 14 67160 54 67480
rect -346 67120 54 67160
rect -346 66760 54 66800
rect -346 66440 -306 66760
rect 14 66440 54 66760
rect -346 66400 54 66440
rect -346 66040 54 66080
rect -346 65720 -306 66040
rect 14 65720 54 66040
rect -346 65680 54 65720
rect -346 65320 54 65360
rect -346 65000 -306 65320
rect 14 65000 54 65320
rect -346 64960 54 65000
rect -346 64600 54 64640
rect -346 64280 -306 64600
rect 14 64280 54 64600
rect -346 64240 54 64280
rect -346 63880 54 63920
rect -346 63560 -306 63880
rect 14 63560 54 63880
rect -346 63520 54 63560
rect -346 63160 54 63200
rect -346 62840 -306 63160
rect 14 62840 54 63160
rect -346 62800 54 62840
rect -346 62440 54 62480
rect -346 62120 -306 62440
rect 14 62120 54 62440
rect -346 62080 54 62120
rect -346 61720 54 61760
rect -346 61400 -306 61720
rect 14 61400 54 61720
rect -346 61360 54 61400
rect -346 61000 54 61040
rect -346 60680 -306 61000
rect 14 60680 54 61000
rect -346 60640 54 60680
rect -346 60280 54 60320
rect -346 59960 -306 60280
rect 14 59960 54 60280
rect -346 59920 54 59960
rect -346 59560 54 59600
rect -346 59240 -306 59560
rect 14 59240 54 59560
rect -346 59200 54 59240
rect -346 58840 54 58880
rect -346 58520 -306 58840
rect 14 58520 54 58840
rect -346 58480 54 58520
rect -346 58120 54 58160
rect -346 57800 -306 58120
rect 14 57800 54 58120
rect -346 57760 54 57800
rect -346 57400 54 57440
rect -346 57080 -306 57400
rect 14 57080 54 57400
rect -346 57040 54 57080
rect -346 56680 54 56720
rect -346 56360 -306 56680
rect 14 56360 54 56680
rect -346 56320 54 56360
rect -346 55960 54 56000
rect -346 55640 -306 55960
rect 14 55640 54 55960
rect -346 55600 54 55640
rect -346 55240 54 55280
rect -346 54920 -306 55240
rect 14 54920 54 55240
rect -346 54880 54 54920
rect -346 54520 54 54560
rect -346 54200 -306 54520
rect 14 54200 54 54520
rect -346 54160 54 54200
rect -346 53800 54 53840
rect -346 53480 -306 53800
rect 14 53480 54 53800
rect -346 53440 54 53480
rect -346 53080 54 53120
rect -346 52760 -306 53080
rect 14 52760 54 53080
rect -346 52720 54 52760
rect -346 52360 54 52400
rect -346 52040 -306 52360
rect 14 52040 54 52360
rect -346 52000 54 52040
rect -346 51640 54 51680
rect -346 51320 -306 51640
rect 14 51320 54 51640
rect -346 51280 54 51320
rect -346 50920 54 50960
rect -346 50600 -306 50920
rect 14 50600 54 50920
rect -346 50560 54 50600
rect -346 50200 54 50240
rect -346 49880 -306 50200
rect 14 49880 54 50200
rect -346 49840 54 49880
rect -346 49480 54 49520
rect -346 49160 -306 49480
rect 14 49160 54 49480
rect -346 49120 54 49160
rect -346 48760 54 48800
rect -346 48440 -306 48760
rect 14 48440 54 48760
rect -346 48400 54 48440
rect -346 48040 54 48080
rect -346 47720 -306 48040
rect 14 47720 54 48040
rect -346 47680 54 47720
rect -346 47320 54 47360
rect -346 47000 -306 47320
rect 14 47000 54 47320
rect -346 46960 54 47000
rect -346 46600 54 46640
rect -346 46280 -306 46600
rect 14 46280 54 46600
rect -346 46240 54 46280
rect -346 45880 54 45920
rect -346 45560 -306 45880
rect 14 45560 54 45880
rect -346 45520 54 45560
rect -346 45160 54 45200
rect -346 44840 -306 45160
rect 14 44840 54 45160
rect -346 44800 54 44840
rect -346 44440 54 44480
rect -346 44120 -306 44440
rect 14 44120 54 44440
rect -346 44080 54 44120
rect -346 43720 54 43760
rect -346 43400 -306 43720
rect 14 43400 54 43720
rect -346 43360 54 43400
rect -346 43000 54 43040
rect -346 42680 -306 43000
rect 14 42680 54 43000
rect -346 42640 54 42680
rect -346 42280 54 42320
rect -346 41960 -306 42280
rect 14 41960 54 42280
rect -346 41920 54 41960
rect -346 41560 54 41600
rect -346 41240 -306 41560
rect 14 41240 54 41560
rect -346 41200 54 41240
rect -346 40840 54 40880
rect -346 40520 -306 40840
rect 14 40520 54 40840
rect -346 40480 54 40520
rect -346 40120 54 40160
rect -346 39800 -306 40120
rect 14 39800 54 40120
rect -346 39760 54 39800
rect -346 39400 54 39440
rect -346 39080 -306 39400
rect 14 39080 54 39400
rect -346 39040 54 39080
rect -346 38680 54 38720
rect -346 38360 -306 38680
rect 14 38360 54 38680
rect -346 38320 54 38360
rect -346 37960 54 38000
rect -346 37640 -306 37960
rect 14 37640 54 37960
rect -346 37600 54 37640
rect -346 37240 54 37280
rect -346 36920 -306 37240
rect 14 36920 54 37240
rect -346 36880 54 36920
rect -346 36520 54 36560
rect -346 36200 -306 36520
rect 14 36200 54 36520
rect -346 36160 54 36200
rect -346 35800 54 35840
rect -346 35480 -306 35800
rect 14 35480 54 35800
rect -346 35440 54 35480
rect -346 35080 54 35120
rect -346 34760 -306 35080
rect 14 34760 54 35080
rect -346 34720 54 34760
rect -346 34360 54 34400
rect -346 34040 -306 34360
rect 14 34040 54 34360
rect -346 34000 54 34040
rect -346 33640 54 33680
rect -346 33320 -306 33640
rect 14 33320 54 33640
rect -346 33280 54 33320
rect -346 32920 54 32960
rect -346 32600 -306 32920
rect 14 32600 54 32920
rect -346 32560 54 32600
rect -346 32200 54 32240
rect -346 31880 -306 32200
rect 14 31880 54 32200
rect -346 31840 54 31880
rect -346 31480 54 31520
rect -346 31160 -306 31480
rect 14 31160 54 31480
rect -346 31120 54 31160
rect -346 30760 54 30800
rect -346 30440 -306 30760
rect 14 30440 54 30760
rect -346 30400 54 30440
rect -346 30040 54 30080
rect -346 29720 -306 30040
rect 14 29720 54 30040
rect -346 29680 54 29720
rect -346 29320 54 29360
rect -346 29000 -306 29320
rect 14 29000 54 29320
rect -346 28960 54 29000
rect -346 28600 54 28640
rect -346 28280 -306 28600
rect 14 28280 54 28600
rect -346 28240 54 28280
rect -346 27880 54 27920
rect -346 27560 -306 27880
rect 14 27560 54 27880
rect -346 27520 54 27560
rect -346 27160 54 27200
rect -346 26840 -306 27160
rect 14 26840 54 27160
rect -346 26800 54 26840
rect -346 26440 54 26480
rect -346 26120 -306 26440
rect 14 26120 54 26440
rect -346 26080 54 26120
rect -346 25720 54 25760
rect -346 25400 -306 25720
rect 14 25400 54 25720
rect -346 25360 54 25400
rect -346 25000 54 25040
rect -346 24680 -306 25000
rect 14 24680 54 25000
rect -346 24640 54 24680
rect -346 24280 54 24320
rect -346 23960 -306 24280
rect 14 23960 54 24280
rect -346 23920 54 23960
rect -346 23560 54 23600
rect -346 23240 -306 23560
rect 14 23240 54 23560
rect -346 23200 54 23240
rect -346 22840 54 22880
rect -346 22520 -306 22840
rect 14 22520 54 22840
rect -346 22480 54 22520
rect -346 22120 54 22160
rect -346 21800 -306 22120
rect 14 21800 54 22120
rect -346 21760 54 21800
rect -346 21400 54 21440
rect -346 21080 -306 21400
rect 14 21080 54 21400
rect -346 21040 54 21080
rect -346 20680 54 20720
rect -346 20360 -306 20680
rect 14 20360 54 20680
rect -346 20320 54 20360
rect -346 19960 54 20000
rect -346 19640 -306 19960
rect 14 19640 54 19960
rect -346 19600 54 19640
rect -346 19240 54 19280
rect -346 18920 -306 19240
rect 14 18920 54 19240
rect -346 18880 54 18920
rect -346 18520 54 18560
rect -346 18200 -306 18520
rect 14 18200 54 18520
rect -346 18160 54 18200
rect -346 17800 54 17840
rect -346 17480 -306 17800
rect 14 17480 54 17800
rect -346 17440 54 17480
rect -346 17080 54 17120
rect -346 16760 -306 17080
rect 14 16760 54 17080
rect -346 16720 54 16760
rect -346 16360 54 16400
rect -346 16040 -306 16360
rect 14 16040 54 16360
rect -346 16000 54 16040
rect -346 15640 54 15680
rect -346 15320 -306 15640
rect 14 15320 54 15640
rect -346 15280 54 15320
rect -346 14920 54 14960
rect -346 14600 -306 14920
rect 14 14600 54 14920
rect -346 14560 54 14600
rect -346 14200 54 14240
rect -346 13880 -306 14200
rect 14 13880 54 14200
rect -346 13840 54 13880
rect -346 13480 54 13520
rect -346 13160 -306 13480
rect 14 13160 54 13480
rect -346 13120 54 13160
rect -346 12760 54 12800
rect -346 12440 -306 12760
rect 14 12440 54 12760
rect -346 12400 54 12440
rect -346 12040 54 12080
rect -346 11720 -306 12040
rect 14 11720 54 12040
rect -346 11680 54 11720
rect -346 11320 54 11360
rect -346 11000 -306 11320
rect 14 11000 54 11320
rect -346 10960 54 11000
rect -346 10600 54 10640
rect -346 10280 -306 10600
rect 14 10280 54 10600
rect -346 10240 54 10280
rect -346 9880 54 9920
rect -346 9560 -306 9880
rect 14 9560 54 9880
rect -346 9520 54 9560
rect -346 9160 54 9200
rect -346 8840 -306 9160
rect 14 8840 54 9160
rect -346 8800 54 8840
rect -346 8440 54 8480
rect -346 8120 -306 8440
rect 14 8120 54 8440
rect -346 8080 54 8120
rect -346 7720 54 7760
rect -346 7400 -306 7720
rect 14 7400 54 7720
rect -346 7360 54 7400
rect -346 7000 54 7040
rect -346 6680 -306 7000
rect 14 6680 54 7000
rect -346 6640 54 6680
rect -346 6280 54 6320
rect -346 5960 -306 6280
rect 14 5960 54 6280
rect -346 5920 54 5960
rect -346 5560 54 5600
rect -346 5240 -306 5560
rect 14 5240 54 5560
rect -346 5200 54 5240
rect -346 4840 54 4880
rect -346 4520 -306 4840
rect 14 4520 54 4840
rect -346 4480 54 4520
rect -346 4120 54 4160
rect -346 3800 -306 4120
rect 14 3800 54 4120
rect -346 3760 54 3800
rect -346 3400 54 3440
rect -346 3080 -306 3400
rect 14 3080 54 3400
rect -346 3040 54 3080
rect -346 2680 54 2720
rect -346 2360 -306 2680
rect 14 2360 54 2680
rect -346 2320 54 2360
rect -346 1960 54 2000
rect -346 1640 -306 1960
rect 14 1640 54 1960
rect -346 1600 54 1640
rect -346 1240 54 1280
rect -346 920 -306 1240
rect 14 920 54 1240
rect -346 880 54 920
rect -346 520 54 560
rect -346 200 -306 520
rect 14 200 54 520
rect -346 160 54 200
rect -346 -200 54 -160
rect -346 -520 -306 -200
rect 14 -520 54 -200
rect -346 -560 54 -520
rect -346 -920 54 -880
rect -346 -1240 -306 -920
rect 14 -1240 54 -920
rect -346 -1280 54 -1240
rect -346 -1640 54 -1600
rect -346 -1960 -306 -1640
rect 14 -1960 54 -1640
rect -346 -2000 54 -1960
rect -346 -2360 54 -2320
rect -346 -2680 -306 -2360
rect 14 -2680 54 -2360
rect -346 -2720 54 -2680
rect -346 -3080 54 -3040
rect -346 -3400 -306 -3080
rect 14 -3400 54 -3080
rect -346 -3440 54 -3400
rect -346 -3800 54 -3760
rect -346 -4120 -306 -3800
rect 14 -4120 54 -3800
rect -346 -4160 54 -4120
rect -346 -4520 54 -4480
rect -346 -4840 -306 -4520
rect 14 -4840 54 -4520
rect -346 -4880 54 -4840
rect -346 -5240 54 -5200
rect -346 -5560 -306 -5240
rect 14 -5560 54 -5240
rect -346 -5600 54 -5560
rect -346 -5960 54 -5920
rect -346 -6280 -306 -5960
rect 14 -6280 54 -5960
rect -346 -6320 54 -6280
rect -346 -6680 54 -6640
rect -346 -7000 -306 -6680
rect 14 -7000 54 -6680
rect -346 -7040 54 -7000
rect -346 -7400 54 -7360
rect -346 -7720 -306 -7400
rect 14 -7720 54 -7400
rect -346 -7760 54 -7720
rect -346 -8120 54 -8080
rect -346 -8440 -306 -8120
rect 14 -8440 54 -8120
rect -346 -8480 54 -8440
rect -346 -8840 54 -8800
rect -346 -9160 -306 -8840
rect 14 -9160 54 -8840
rect -346 -9200 54 -9160
rect -346 -9560 54 -9520
rect -346 -9880 -306 -9560
rect 14 -9880 54 -9560
rect -346 -9920 54 -9880
rect -346 -10280 54 -10240
rect -346 -10600 -306 -10280
rect 14 -10600 54 -10280
rect -346 -10640 54 -10600
rect -346 -11000 54 -10960
rect -346 -11320 -306 -11000
rect 14 -11320 54 -11000
rect -346 -11360 54 -11320
rect -346 -11720 54 -11680
rect -346 -12040 -306 -11720
rect 14 -12040 54 -11720
rect -346 -12080 54 -12040
rect -346 -12440 54 -12400
rect -346 -12760 -306 -12440
rect 14 -12760 54 -12440
rect -346 -12800 54 -12760
rect -346 -13160 54 -13120
rect -346 -13480 -306 -13160
rect 14 -13480 54 -13160
rect -346 -13520 54 -13480
rect -346 -13880 54 -13840
rect -346 -14200 -306 -13880
rect 14 -14200 54 -13880
rect -346 -14240 54 -14200
rect -346 -14600 54 -14560
rect -346 -14920 -306 -14600
rect 14 -14920 54 -14600
rect -346 -14960 54 -14920
rect -346 -15320 54 -15280
rect -346 -15640 -306 -15320
rect 14 -15640 54 -15320
rect -346 -15680 54 -15640
rect -346 -16040 54 -16000
rect -346 -16360 -306 -16040
rect 14 -16360 54 -16040
rect -346 -16400 54 -16360
rect -346 -16760 54 -16720
rect -346 -17080 -306 -16760
rect 14 -17080 54 -16760
rect -346 -17120 54 -17080
rect -346 -17480 54 -17440
rect -346 -17800 -306 -17480
rect 14 -17800 54 -17480
rect -346 -17840 54 -17800
rect -346 -18200 54 -18160
rect -346 -18520 -306 -18200
rect 14 -18520 54 -18200
rect -346 -18560 54 -18520
rect -346 -18920 54 -18880
rect -346 -19240 -306 -18920
rect 14 -19240 54 -18920
rect -346 -19280 54 -19240
rect -346 -19640 54 -19600
rect -346 -19960 -306 -19640
rect 14 -19960 54 -19640
rect -346 -20000 54 -19960
rect -346 -20360 54 -20320
rect -346 -20680 -306 -20360
rect 14 -20680 54 -20360
rect -346 -20720 54 -20680
rect -346 -21080 54 -21040
rect -346 -21400 -306 -21080
rect 14 -21400 54 -21080
rect -346 -21440 54 -21400
rect -346 -21800 54 -21760
rect -346 -22120 -306 -21800
rect 14 -22120 54 -21800
rect -346 -22160 54 -22120
rect -346 -22520 54 -22480
rect -346 -22840 -306 -22520
rect 14 -22840 54 -22520
rect -346 -22880 54 -22840
rect -346 -23240 54 -23200
rect -346 -23560 -306 -23240
rect 14 -23560 54 -23240
rect -346 -23600 54 -23560
rect -346 -23960 54 -23920
rect -346 -24280 -306 -23960
rect 14 -24280 54 -23960
rect -346 -24320 54 -24280
rect -346 -24680 54 -24640
rect -346 -25000 -306 -24680
rect 14 -25000 54 -24680
rect -346 -25040 54 -25000
rect -346 -25400 54 -25360
rect -346 -25720 -306 -25400
rect 14 -25720 54 -25400
rect -346 -25760 54 -25720
rect -346 -26120 54 -26080
rect -346 -26440 -306 -26120
rect 14 -26440 54 -26120
rect -346 -26480 54 -26440
rect -346 -26840 54 -26800
rect -346 -27160 -306 -26840
rect 14 -27160 54 -26840
rect -346 -27200 54 -27160
rect -346 -27560 54 -27520
rect -346 -27880 -306 -27560
rect 14 -27880 54 -27560
rect -346 -27920 54 -27880
rect -346 -28280 54 -28240
rect -346 -28600 -306 -28280
rect 14 -28600 54 -28280
rect -346 -28640 54 -28600
rect -346 -29000 54 -28960
rect -346 -29320 -306 -29000
rect 14 -29320 54 -29000
rect -346 -29360 54 -29320
rect -346 -29720 54 -29680
rect -346 -30040 -306 -29720
rect 14 -30040 54 -29720
rect -346 -30080 54 -30040
rect -346 -30440 54 -30400
rect -346 -30760 -306 -30440
rect 14 -30760 54 -30440
rect -346 -30800 54 -30760
rect -346 -31160 54 -31120
rect -346 -31480 -306 -31160
rect 14 -31480 54 -31160
rect -346 -31520 54 -31480
rect -346 -31880 54 -31840
rect -346 -32200 -306 -31880
rect 14 -32200 54 -31880
rect -346 -32240 54 -32200
rect -346 -32600 54 -32560
rect -346 -32920 -306 -32600
rect 14 -32920 54 -32600
rect -346 -32960 54 -32920
rect -346 -33320 54 -33280
rect -346 -33640 -306 -33320
rect 14 -33640 54 -33320
rect -346 -33680 54 -33640
rect -346 -34040 54 -34000
rect -346 -34360 -306 -34040
rect 14 -34360 54 -34040
rect -346 -34400 54 -34360
rect -346 -34760 54 -34720
rect -346 -35080 -306 -34760
rect 14 -35080 54 -34760
rect -346 -35120 54 -35080
rect -346 -35480 54 -35440
rect -346 -35800 -306 -35480
rect 14 -35800 54 -35480
rect -346 -35840 54 -35800
rect -346 -36200 54 -36160
rect -346 -36520 -306 -36200
rect 14 -36520 54 -36200
rect -346 -36560 54 -36520
rect -346 -36920 54 -36880
rect -346 -37240 -306 -36920
rect 14 -37240 54 -36920
rect -346 -37280 54 -37240
rect -346 -37640 54 -37600
rect -346 -37960 -306 -37640
rect 14 -37960 54 -37640
rect -346 -38000 54 -37960
rect -346 -38360 54 -38320
rect -346 -38680 -306 -38360
rect 14 -38680 54 -38360
rect -346 -38720 54 -38680
rect -346 -39080 54 -39040
rect -346 -39400 -306 -39080
rect 14 -39400 54 -39080
rect -346 -39440 54 -39400
rect -346 -39800 54 -39760
rect -346 -40120 -306 -39800
rect 14 -40120 54 -39800
rect -346 -40160 54 -40120
rect -346 -40520 54 -40480
rect -346 -40840 -306 -40520
rect 14 -40840 54 -40520
rect -346 -40880 54 -40840
rect -346 -41240 54 -41200
rect -346 -41560 -306 -41240
rect 14 -41560 54 -41240
rect -346 -41600 54 -41560
rect -346 -41960 54 -41920
rect -346 -42280 -306 -41960
rect 14 -42280 54 -41960
rect -346 -42320 54 -42280
rect -346 -42680 54 -42640
rect -346 -43000 -306 -42680
rect 14 -43000 54 -42680
rect -346 -43040 54 -43000
rect -346 -43400 54 -43360
rect -346 -43720 -306 -43400
rect 14 -43720 54 -43400
rect -346 -43760 54 -43720
rect -346 -44120 54 -44080
rect -346 -44440 -306 -44120
rect 14 -44440 54 -44120
rect -346 -44480 54 -44440
rect -346 -44840 54 -44800
rect -346 -45160 -306 -44840
rect 14 -45160 54 -44840
rect -346 -45200 54 -45160
rect -346 -45560 54 -45520
rect -346 -45880 -306 -45560
rect 14 -45880 54 -45560
rect -346 -45920 54 -45880
rect -346 -46280 54 -46240
rect -346 -46600 -306 -46280
rect 14 -46600 54 -46280
rect -346 -46640 54 -46600
rect -346 -47000 54 -46960
rect -346 -47320 -306 -47000
rect 14 -47320 54 -47000
rect -346 -47360 54 -47320
rect -346 -47720 54 -47680
rect -346 -48040 -306 -47720
rect 14 -48040 54 -47720
rect -346 -48080 54 -48040
rect -346 -48440 54 -48400
rect -346 -48760 -306 -48440
rect 14 -48760 54 -48440
rect -346 -48800 54 -48760
rect -346 -49160 54 -49120
rect -346 -49480 -306 -49160
rect 14 -49480 54 -49160
rect -346 -49520 54 -49480
rect -346 -49880 54 -49840
rect -346 -50200 -306 -49880
rect 14 -50200 54 -49880
rect -346 -50240 54 -50200
rect -346 -50600 54 -50560
rect -346 -50920 -306 -50600
rect 14 -50920 54 -50600
rect -346 -50960 54 -50920
rect -346 -51320 54 -51280
rect -346 -51640 -306 -51320
rect 14 -51640 54 -51320
rect -346 -51680 54 -51640
rect -346 -52040 54 -52000
rect -346 -52360 -306 -52040
rect 14 -52360 54 -52040
rect -346 -52400 54 -52360
rect -346 -52760 54 -52720
rect -346 -53080 -306 -52760
rect 14 -53080 54 -52760
rect -346 -53120 54 -53080
rect -346 -53480 54 -53440
rect -346 -53800 -306 -53480
rect 14 -53800 54 -53480
rect -346 -53840 54 -53800
rect -346 -54200 54 -54160
rect -346 -54520 -306 -54200
rect 14 -54520 54 -54200
rect -346 -54560 54 -54520
rect -346 -54920 54 -54880
rect -346 -55240 -306 -54920
rect 14 -55240 54 -54920
rect -346 -55280 54 -55240
rect -346 -55640 54 -55600
rect -346 -55960 -306 -55640
rect 14 -55960 54 -55640
rect -346 -56000 54 -55960
rect -346 -56360 54 -56320
rect -346 -56680 -306 -56360
rect 14 -56680 54 -56360
rect -346 -56720 54 -56680
rect -346 -57080 54 -57040
rect -346 -57400 -306 -57080
rect 14 -57400 54 -57080
rect -346 -57440 54 -57400
rect -346 -57800 54 -57760
rect -346 -58120 -306 -57800
rect 14 -58120 54 -57800
rect -346 -58160 54 -58120
rect -346 -58520 54 -58480
rect -346 -58840 -306 -58520
rect 14 -58840 54 -58520
rect -346 -58880 54 -58840
rect -346 -59240 54 -59200
rect -346 -59560 -306 -59240
rect 14 -59560 54 -59240
rect -346 -59600 54 -59560
rect -346 -59960 54 -59920
rect -346 -60280 -306 -59960
rect 14 -60280 54 -59960
rect -346 -60320 54 -60280
rect -346 -60680 54 -60640
rect -346 -61000 -306 -60680
rect 14 -61000 54 -60680
rect -346 -61040 54 -61000
rect -346 -61400 54 -61360
rect -346 -61720 -306 -61400
rect 14 -61720 54 -61400
rect -346 -61760 54 -61720
rect -346 -62120 54 -62080
rect -346 -62440 -306 -62120
rect 14 -62440 54 -62120
rect -346 -62480 54 -62440
rect -346 -62840 54 -62800
rect -346 -63160 -306 -62840
rect 14 -63160 54 -62840
rect -346 -63200 54 -63160
rect -346 -63560 54 -63520
rect -346 -63880 -306 -63560
rect 14 -63880 54 -63560
rect -346 -63920 54 -63880
rect -346 -64280 54 -64240
rect -346 -64600 -306 -64280
rect 14 -64600 54 -64280
rect -346 -64640 54 -64600
rect -346 -65000 54 -64960
rect -346 -65320 -306 -65000
rect 14 -65320 54 -65000
rect -346 -65360 54 -65320
rect -346 -65720 54 -65680
rect -346 -66040 -306 -65720
rect 14 -66040 54 -65720
rect -346 -66080 54 -66040
rect -346 -66440 54 -66400
rect -346 -66760 -306 -66440
rect 14 -66760 54 -66440
rect -346 -66800 54 -66760
rect -346 -67160 54 -67120
rect -346 -67480 -306 -67160
rect 14 -67480 54 -67160
rect -346 -67520 54 -67480
rect -346 -67880 54 -67840
rect -346 -68200 -306 -67880
rect 14 -68200 54 -67880
rect -346 -68240 54 -68200
rect -346 -68600 54 -68560
rect -346 -68920 -306 -68600
rect 14 -68920 54 -68600
rect -346 -68960 54 -68920
rect -346 -69320 54 -69280
rect -346 -69640 -306 -69320
rect 14 -69640 54 -69320
rect -346 -69680 54 -69640
rect -346 -70040 54 -70000
rect -346 -70360 -306 -70040
rect 14 -70360 54 -70040
rect -346 -70400 54 -70360
rect -346 -70760 54 -70720
rect -346 -71080 -306 -70760
rect 14 -71080 54 -70760
rect -346 -71120 54 -71080
rect -346 -71480 54 -71440
rect -346 -71800 -306 -71480
rect 14 -71800 54 -71480
rect -346 -71840 54 -71800
rect -346 -72200 54 -72160
rect -346 -72520 -306 -72200
rect 14 -72520 54 -72200
rect -346 -72560 54 -72520
rect -346 -72920 54 -72880
rect -346 -73240 -306 -72920
rect 14 -73240 54 -72920
rect -346 -73280 54 -73240
rect -346 -73640 54 -73600
rect -346 -73960 -306 -73640
rect 14 -73960 54 -73640
rect -346 -74000 54 -73960
rect -346 -74360 54 -74320
rect -346 -74680 -306 -74360
rect 14 -74680 54 -74360
rect -346 -74720 54 -74680
rect -346 -75080 54 -75040
rect -346 -75400 -306 -75080
rect 14 -75400 54 -75080
rect -346 -75440 54 -75400
rect -346 -75800 54 -75760
rect -346 -76120 -306 -75800
rect 14 -76120 54 -75800
rect -346 -76160 54 -76120
rect -346 -76520 54 -76480
rect -346 -76840 -306 -76520
rect 14 -76840 54 -76520
rect -346 -76880 54 -76840
rect -346 -77240 54 -77200
rect -346 -77560 -306 -77240
rect 14 -77560 54 -77240
rect -346 -77600 54 -77560
rect -346 -77960 54 -77920
rect -346 -78280 -306 -77960
rect 14 -78280 54 -77960
rect -346 -78320 54 -78280
rect -346 -78680 54 -78640
rect -346 -79000 -306 -78680
rect 14 -79000 54 -78680
rect -346 -79040 54 -79000
rect -346 -79400 54 -79360
rect -346 -79720 -306 -79400
rect 14 -79720 54 -79400
rect -346 -79760 54 -79720
rect -346 -80120 54 -80080
rect -346 -80440 -306 -80120
rect 14 -80440 54 -80120
rect -346 -80480 54 -80440
rect -346 -80840 54 -80800
rect -346 -81160 -306 -80840
rect 14 -81160 54 -80840
rect -346 -81200 54 -81160
rect -346 -81560 54 -81520
rect -346 -81880 -306 -81560
rect 14 -81880 54 -81560
rect -346 -81920 54 -81880
rect -346 -82280 54 -82240
rect -346 -82600 -306 -82280
rect 14 -82600 54 -82280
rect -346 -82640 54 -82600
rect -346 -83000 54 -82960
rect -346 -83320 -306 -83000
rect 14 -83320 54 -83000
rect -346 -83360 54 -83320
rect -346 -83720 54 -83680
rect -346 -84040 -306 -83720
rect 14 -84040 54 -83720
rect -346 -84080 54 -84040
rect -346 -84440 54 -84400
rect -346 -84760 -306 -84440
rect 14 -84760 54 -84440
rect -346 -84800 54 -84760
rect -346 -85160 54 -85120
rect -346 -85480 -306 -85160
rect 14 -85480 54 -85160
rect -346 -85520 54 -85480
rect -346 -85880 54 -85840
rect -346 -86200 -306 -85880
rect 14 -86200 54 -85880
rect -346 -86240 54 -86200
rect -346 -86600 54 -86560
rect -346 -86920 -306 -86600
rect 14 -86920 54 -86600
rect -346 -86960 54 -86920
rect -346 -87320 54 -87280
rect -346 -87640 -306 -87320
rect 14 -87640 54 -87320
rect -346 -87680 54 -87640
rect -346 -88040 54 -88000
rect -346 -88360 -306 -88040
rect 14 -88360 54 -88040
rect -346 -88400 54 -88360
rect -346 -88760 54 -88720
rect -346 -89080 -306 -88760
rect 14 -89080 54 -88760
rect -346 -89120 54 -89080
rect -346 -89480 54 -89440
rect -346 -89800 -306 -89480
rect 14 -89800 54 -89480
rect -346 -89840 54 -89800
rect -346 -90200 54 -90160
rect -346 -90520 -306 -90200
rect 14 -90520 54 -90200
rect -346 -90560 54 -90520
rect -346 -90920 54 -90880
rect -346 -91240 -306 -90920
rect 14 -91240 54 -90920
rect -346 -91280 54 -91240
rect -346 -91640 54 -91600
rect -346 -91960 -306 -91640
rect 14 -91960 54 -91640
rect -346 -92000 54 -91960
<< mimcapcontact >>
rect -306 91640 14 91960
rect -306 90920 14 91240
rect -306 90200 14 90520
rect -306 89480 14 89800
rect -306 88760 14 89080
rect -306 88040 14 88360
rect -306 87320 14 87640
rect -306 86600 14 86920
rect -306 85880 14 86200
rect -306 85160 14 85480
rect -306 84440 14 84760
rect -306 83720 14 84040
rect -306 83000 14 83320
rect -306 82280 14 82600
rect -306 81560 14 81880
rect -306 80840 14 81160
rect -306 80120 14 80440
rect -306 79400 14 79720
rect -306 78680 14 79000
rect -306 77960 14 78280
rect -306 77240 14 77560
rect -306 76520 14 76840
rect -306 75800 14 76120
rect -306 75080 14 75400
rect -306 74360 14 74680
rect -306 73640 14 73960
rect -306 72920 14 73240
rect -306 72200 14 72520
rect -306 71480 14 71800
rect -306 70760 14 71080
rect -306 70040 14 70360
rect -306 69320 14 69640
rect -306 68600 14 68920
rect -306 67880 14 68200
rect -306 67160 14 67480
rect -306 66440 14 66760
rect -306 65720 14 66040
rect -306 65000 14 65320
rect -306 64280 14 64600
rect -306 63560 14 63880
rect -306 62840 14 63160
rect -306 62120 14 62440
rect -306 61400 14 61720
rect -306 60680 14 61000
rect -306 59960 14 60280
rect -306 59240 14 59560
rect -306 58520 14 58840
rect -306 57800 14 58120
rect -306 57080 14 57400
rect -306 56360 14 56680
rect -306 55640 14 55960
rect -306 54920 14 55240
rect -306 54200 14 54520
rect -306 53480 14 53800
rect -306 52760 14 53080
rect -306 52040 14 52360
rect -306 51320 14 51640
rect -306 50600 14 50920
rect -306 49880 14 50200
rect -306 49160 14 49480
rect -306 48440 14 48760
rect -306 47720 14 48040
rect -306 47000 14 47320
rect -306 46280 14 46600
rect -306 45560 14 45880
rect -306 44840 14 45160
rect -306 44120 14 44440
rect -306 43400 14 43720
rect -306 42680 14 43000
rect -306 41960 14 42280
rect -306 41240 14 41560
rect -306 40520 14 40840
rect -306 39800 14 40120
rect -306 39080 14 39400
rect -306 38360 14 38680
rect -306 37640 14 37960
rect -306 36920 14 37240
rect -306 36200 14 36520
rect -306 35480 14 35800
rect -306 34760 14 35080
rect -306 34040 14 34360
rect -306 33320 14 33640
rect -306 32600 14 32920
rect -306 31880 14 32200
rect -306 31160 14 31480
rect -306 30440 14 30760
rect -306 29720 14 30040
rect -306 29000 14 29320
rect -306 28280 14 28600
rect -306 27560 14 27880
rect -306 26840 14 27160
rect -306 26120 14 26440
rect -306 25400 14 25720
rect -306 24680 14 25000
rect -306 23960 14 24280
rect -306 23240 14 23560
rect -306 22520 14 22840
rect -306 21800 14 22120
rect -306 21080 14 21400
rect -306 20360 14 20680
rect -306 19640 14 19960
rect -306 18920 14 19240
rect -306 18200 14 18520
rect -306 17480 14 17800
rect -306 16760 14 17080
rect -306 16040 14 16360
rect -306 15320 14 15640
rect -306 14600 14 14920
rect -306 13880 14 14200
rect -306 13160 14 13480
rect -306 12440 14 12760
rect -306 11720 14 12040
rect -306 11000 14 11320
rect -306 10280 14 10600
rect -306 9560 14 9880
rect -306 8840 14 9160
rect -306 8120 14 8440
rect -306 7400 14 7720
rect -306 6680 14 7000
rect -306 5960 14 6280
rect -306 5240 14 5560
rect -306 4520 14 4840
rect -306 3800 14 4120
rect -306 3080 14 3400
rect -306 2360 14 2680
rect -306 1640 14 1960
rect -306 920 14 1240
rect -306 200 14 520
rect -306 -520 14 -200
rect -306 -1240 14 -920
rect -306 -1960 14 -1640
rect -306 -2680 14 -2360
rect -306 -3400 14 -3080
rect -306 -4120 14 -3800
rect -306 -4840 14 -4520
rect -306 -5560 14 -5240
rect -306 -6280 14 -5960
rect -306 -7000 14 -6680
rect -306 -7720 14 -7400
rect -306 -8440 14 -8120
rect -306 -9160 14 -8840
rect -306 -9880 14 -9560
rect -306 -10600 14 -10280
rect -306 -11320 14 -11000
rect -306 -12040 14 -11720
rect -306 -12760 14 -12440
rect -306 -13480 14 -13160
rect -306 -14200 14 -13880
rect -306 -14920 14 -14600
rect -306 -15640 14 -15320
rect -306 -16360 14 -16040
rect -306 -17080 14 -16760
rect -306 -17800 14 -17480
rect -306 -18520 14 -18200
rect -306 -19240 14 -18920
rect -306 -19960 14 -19640
rect -306 -20680 14 -20360
rect -306 -21400 14 -21080
rect -306 -22120 14 -21800
rect -306 -22840 14 -22520
rect -306 -23560 14 -23240
rect -306 -24280 14 -23960
rect -306 -25000 14 -24680
rect -306 -25720 14 -25400
rect -306 -26440 14 -26120
rect -306 -27160 14 -26840
rect -306 -27880 14 -27560
rect -306 -28600 14 -28280
rect -306 -29320 14 -29000
rect -306 -30040 14 -29720
rect -306 -30760 14 -30440
rect -306 -31480 14 -31160
rect -306 -32200 14 -31880
rect -306 -32920 14 -32600
rect -306 -33640 14 -33320
rect -306 -34360 14 -34040
rect -306 -35080 14 -34760
rect -306 -35800 14 -35480
rect -306 -36520 14 -36200
rect -306 -37240 14 -36920
rect -306 -37960 14 -37640
rect -306 -38680 14 -38360
rect -306 -39400 14 -39080
rect -306 -40120 14 -39800
rect -306 -40840 14 -40520
rect -306 -41560 14 -41240
rect -306 -42280 14 -41960
rect -306 -43000 14 -42680
rect -306 -43720 14 -43400
rect -306 -44440 14 -44120
rect -306 -45160 14 -44840
rect -306 -45880 14 -45560
rect -306 -46600 14 -46280
rect -306 -47320 14 -47000
rect -306 -48040 14 -47720
rect -306 -48760 14 -48440
rect -306 -49480 14 -49160
rect -306 -50200 14 -49880
rect -306 -50920 14 -50600
rect -306 -51640 14 -51320
rect -306 -52360 14 -52040
rect -306 -53080 14 -52760
rect -306 -53800 14 -53480
rect -306 -54520 14 -54200
rect -306 -55240 14 -54920
rect -306 -55960 14 -55640
rect -306 -56680 14 -56360
rect -306 -57400 14 -57080
rect -306 -58120 14 -57800
rect -306 -58840 14 -58520
rect -306 -59560 14 -59240
rect -306 -60280 14 -59960
rect -306 -61000 14 -60680
rect -306 -61720 14 -61400
rect -306 -62440 14 -62120
rect -306 -63160 14 -62840
rect -306 -63880 14 -63560
rect -306 -64600 14 -64280
rect -306 -65320 14 -65000
rect -306 -66040 14 -65720
rect -306 -66760 14 -66440
rect -306 -67480 14 -67160
rect -306 -68200 14 -67880
rect -306 -68920 14 -68600
rect -306 -69640 14 -69320
rect -306 -70360 14 -70040
rect -306 -71080 14 -70760
rect -306 -71800 14 -71480
rect -306 -72520 14 -72200
rect -306 -73240 14 -72920
rect -306 -73960 14 -73640
rect -306 -74680 14 -74360
rect -306 -75400 14 -75080
rect -306 -76120 14 -75800
rect -306 -76840 14 -76520
rect -306 -77560 14 -77240
rect -306 -78280 14 -77960
rect -306 -79000 14 -78680
rect -306 -79720 14 -79400
rect -306 -80440 14 -80120
rect -306 -81160 14 -80840
rect -306 -81880 14 -81560
rect -306 -82600 14 -82280
rect -306 -83320 14 -83000
rect -306 -84040 14 -83720
rect -306 -84760 14 -84440
rect -306 -85480 14 -85160
rect -306 -86200 14 -85880
rect -306 -86920 14 -86600
rect -306 -87640 14 -87320
rect -306 -88360 14 -88040
rect -306 -89080 14 -88760
rect -306 -89800 14 -89480
rect -306 -90520 14 -90200
rect -306 -91240 14 -90920
rect -306 -91960 14 -91640
<< metal4 >>
rect -198 91961 -94 92160
rect 282 92012 386 92160
rect -307 91960 15 91961
rect -307 91640 -306 91960
rect 14 91640 15 91960
rect -307 91639 15 91640
rect -198 91241 -94 91639
rect 282 91588 302 92012
rect 366 91588 386 92012
rect 282 91292 386 91588
rect -307 91240 15 91241
rect -307 90920 -306 91240
rect 14 90920 15 91240
rect -307 90919 15 90920
rect -198 90521 -94 90919
rect 282 90868 302 91292
rect 366 90868 386 91292
rect 282 90572 386 90868
rect -307 90520 15 90521
rect -307 90200 -306 90520
rect 14 90200 15 90520
rect -307 90199 15 90200
rect -198 89801 -94 90199
rect 282 90148 302 90572
rect 366 90148 386 90572
rect 282 89852 386 90148
rect -307 89800 15 89801
rect -307 89480 -306 89800
rect 14 89480 15 89800
rect -307 89479 15 89480
rect -198 89081 -94 89479
rect 282 89428 302 89852
rect 366 89428 386 89852
rect 282 89132 386 89428
rect -307 89080 15 89081
rect -307 88760 -306 89080
rect 14 88760 15 89080
rect -307 88759 15 88760
rect -198 88361 -94 88759
rect 282 88708 302 89132
rect 366 88708 386 89132
rect 282 88412 386 88708
rect -307 88360 15 88361
rect -307 88040 -306 88360
rect 14 88040 15 88360
rect -307 88039 15 88040
rect -198 87641 -94 88039
rect 282 87988 302 88412
rect 366 87988 386 88412
rect 282 87692 386 87988
rect -307 87640 15 87641
rect -307 87320 -306 87640
rect 14 87320 15 87640
rect -307 87319 15 87320
rect -198 86921 -94 87319
rect 282 87268 302 87692
rect 366 87268 386 87692
rect 282 86972 386 87268
rect -307 86920 15 86921
rect -307 86600 -306 86920
rect 14 86600 15 86920
rect -307 86599 15 86600
rect -198 86201 -94 86599
rect 282 86548 302 86972
rect 366 86548 386 86972
rect 282 86252 386 86548
rect -307 86200 15 86201
rect -307 85880 -306 86200
rect 14 85880 15 86200
rect -307 85879 15 85880
rect -198 85481 -94 85879
rect 282 85828 302 86252
rect 366 85828 386 86252
rect 282 85532 386 85828
rect -307 85480 15 85481
rect -307 85160 -306 85480
rect 14 85160 15 85480
rect -307 85159 15 85160
rect -198 84761 -94 85159
rect 282 85108 302 85532
rect 366 85108 386 85532
rect 282 84812 386 85108
rect -307 84760 15 84761
rect -307 84440 -306 84760
rect 14 84440 15 84760
rect -307 84439 15 84440
rect -198 84041 -94 84439
rect 282 84388 302 84812
rect 366 84388 386 84812
rect 282 84092 386 84388
rect -307 84040 15 84041
rect -307 83720 -306 84040
rect 14 83720 15 84040
rect -307 83719 15 83720
rect -198 83321 -94 83719
rect 282 83668 302 84092
rect 366 83668 386 84092
rect 282 83372 386 83668
rect -307 83320 15 83321
rect -307 83000 -306 83320
rect 14 83000 15 83320
rect -307 82999 15 83000
rect -198 82601 -94 82999
rect 282 82948 302 83372
rect 366 82948 386 83372
rect 282 82652 386 82948
rect -307 82600 15 82601
rect -307 82280 -306 82600
rect 14 82280 15 82600
rect -307 82279 15 82280
rect -198 81881 -94 82279
rect 282 82228 302 82652
rect 366 82228 386 82652
rect 282 81932 386 82228
rect -307 81880 15 81881
rect -307 81560 -306 81880
rect 14 81560 15 81880
rect -307 81559 15 81560
rect -198 81161 -94 81559
rect 282 81508 302 81932
rect 366 81508 386 81932
rect 282 81212 386 81508
rect -307 81160 15 81161
rect -307 80840 -306 81160
rect 14 80840 15 81160
rect -307 80839 15 80840
rect -198 80441 -94 80839
rect 282 80788 302 81212
rect 366 80788 386 81212
rect 282 80492 386 80788
rect -307 80440 15 80441
rect -307 80120 -306 80440
rect 14 80120 15 80440
rect -307 80119 15 80120
rect -198 79721 -94 80119
rect 282 80068 302 80492
rect 366 80068 386 80492
rect 282 79772 386 80068
rect -307 79720 15 79721
rect -307 79400 -306 79720
rect 14 79400 15 79720
rect -307 79399 15 79400
rect -198 79001 -94 79399
rect 282 79348 302 79772
rect 366 79348 386 79772
rect 282 79052 386 79348
rect -307 79000 15 79001
rect -307 78680 -306 79000
rect 14 78680 15 79000
rect -307 78679 15 78680
rect -198 78281 -94 78679
rect 282 78628 302 79052
rect 366 78628 386 79052
rect 282 78332 386 78628
rect -307 78280 15 78281
rect -307 77960 -306 78280
rect 14 77960 15 78280
rect -307 77959 15 77960
rect -198 77561 -94 77959
rect 282 77908 302 78332
rect 366 77908 386 78332
rect 282 77612 386 77908
rect -307 77560 15 77561
rect -307 77240 -306 77560
rect 14 77240 15 77560
rect -307 77239 15 77240
rect -198 76841 -94 77239
rect 282 77188 302 77612
rect 366 77188 386 77612
rect 282 76892 386 77188
rect -307 76840 15 76841
rect -307 76520 -306 76840
rect 14 76520 15 76840
rect -307 76519 15 76520
rect -198 76121 -94 76519
rect 282 76468 302 76892
rect 366 76468 386 76892
rect 282 76172 386 76468
rect -307 76120 15 76121
rect -307 75800 -306 76120
rect 14 75800 15 76120
rect -307 75799 15 75800
rect -198 75401 -94 75799
rect 282 75748 302 76172
rect 366 75748 386 76172
rect 282 75452 386 75748
rect -307 75400 15 75401
rect -307 75080 -306 75400
rect 14 75080 15 75400
rect -307 75079 15 75080
rect -198 74681 -94 75079
rect 282 75028 302 75452
rect 366 75028 386 75452
rect 282 74732 386 75028
rect -307 74680 15 74681
rect -307 74360 -306 74680
rect 14 74360 15 74680
rect -307 74359 15 74360
rect -198 73961 -94 74359
rect 282 74308 302 74732
rect 366 74308 386 74732
rect 282 74012 386 74308
rect -307 73960 15 73961
rect -307 73640 -306 73960
rect 14 73640 15 73960
rect -307 73639 15 73640
rect -198 73241 -94 73639
rect 282 73588 302 74012
rect 366 73588 386 74012
rect 282 73292 386 73588
rect -307 73240 15 73241
rect -307 72920 -306 73240
rect 14 72920 15 73240
rect -307 72919 15 72920
rect -198 72521 -94 72919
rect 282 72868 302 73292
rect 366 72868 386 73292
rect 282 72572 386 72868
rect -307 72520 15 72521
rect -307 72200 -306 72520
rect 14 72200 15 72520
rect -307 72199 15 72200
rect -198 71801 -94 72199
rect 282 72148 302 72572
rect 366 72148 386 72572
rect 282 71852 386 72148
rect -307 71800 15 71801
rect -307 71480 -306 71800
rect 14 71480 15 71800
rect -307 71479 15 71480
rect -198 71081 -94 71479
rect 282 71428 302 71852
rect 366 71428 386 71852
rect 282 71132 386 71428
rect -307 71080 15 71081
rect -307 70760 -306 71080
rect 14 70760 15 71080
rect -307 70759 15 70760
rect -198 70361 -94 70759
rect 282 70708 302 71132
rect 366 70708 386 71132
rect 282 70412 386 70708
rect -307 70360 15 70361
rect -307 70040 -306 70360
rect 14 70040 15 70360
rect -307 70039 15 70040
rect -198 69641 -94 70039
rect 282 69988 302 70412
rect 366 69988 386 70412
rect 282 69692 386 69988
rect -307 69640 15 69641
rect -307 69320 -306 69640
rect 14 69320 15 69640
rect -307 69319 15 69320
rect -198 68921 -94 69319
rect 282 69268 302 69692
rect 366 69268 386 69692
rect 282 68972 386 69268
rect -307 68920 15 68921
rect -307 68600 -306 68920
rect 14 68600 15 68920
rect -307 68599 15 68600
rect -198 68201 -94 68599
rect 282 68548 302 68972
rect 366 68548 386 68972
rect 282 68252 386 68548
rect -307 68200 15 68201
rect -307 67880 -306 68200
rect 14 67880 15 68200
rect -307 67879 15 67880
rect -198 67481 -94 67879
rect 282 67828 302 68252
rect 366 67828 386 68252
rect 282 67532 386 67828
rect -307 67480 15 67481
rect -307 67160 -306 67480
rect 14 67160 15 67480
rect -307 67159 15 67160
rect -198 66761 -94 67159
rect 282 67108 302 67532
rect 366 67108 386 67532
rect 282 66812 386 67108
rect -307 66760 15 66761
rect -307 66440 -306 66760
rect 14 66440 15 66760
rect -307 66439 15 66440
rect -198 66041 -94 66439
rect 282 66388 302 66812
rect 366 66388 386 66812
rect 282 66092 386 66388
rect -307 66040 15 66041
rect -307 65720 -306 66040
rect 14 65720 15 66040
rect -307 65719 15 65720
rect -198 65321 -94 65719
rect 282 65668 302 66092
rect 366 65668 386 66092
rect 282 65372 386 65668
rect -307 65320 15 65321
rect -307 65000 -306 65320
rect 14 65000 15 65320
rect -307 64999 15 65000
rect -198 64601 -94 64999
rect 282 64948 302 65372
rect 366 64948 386 65372
rect 282 64652 386 64948
rect -307 64600 15 64601
rect -307 64280 -306 64600
rect 14 64280 15 64600
rect -307 64279 15 64280
rect -198 63881 -94 64279
rect 282 64228 302 64652
rect 366 64228 386 64652
rect 282 63932 386 64228
rect -307 63880 15 63881
rect -307 63560 -306 63880
rect 14 63560 15 63880
rect -307 63559 15 63560
rect -198 63161 -94 63559
rect 282 63508 302 63932
rect 366 63508 386 63932
rect 282 63212 386 63508
rect -307 63160 15 63161
rect -307 62840 -306 63160
rect 14 62840 15 63160
rect -307 62839 15 62840
rect -198 62441 -94 62839
rect 282 62788 302 63212
rect 366 62788 386 63212
rect 282 62492 386 62788
rect -307 62440 15 62441
rect -307 62120 -306 62440
rect 14 62120 15 62440
rect -307 62119 15 62120
rect -198 61721 -94 62119
rect 282 62068 302 62492
rect 366 62068 386 62492
rect 282 61772 386 62068
rect -307 61720 15 61721
rect -307 61400 -306 61720
rect 14 61400 15 61720
rect -307 61399 15 61400
rect -198 61001 -94 61399
rect 282 61348 302 61772
rect 366 61348 386 61772
rect 282 61052 386 61348
rect -307 61000 15 61001
rect -307 60680 -306 61000
rect 14 60680 15 61000
rect -307 60679 15 60680
rect -198 60281 -94 60679
rect 282 60628 302 61052
rect 366 60628 386 61052
rect 282 60332 386 60628
rect -307 60280 15 60281
rect -307 59960 -306 60280
rect 14 59960 15 60280
rect -307 59959 15 59960
rect -198 59561 -94 59959
rect 282 59908 302 60332
rect 366 59908 386 60332
rect 282 59612 386 59908
rect -307 59560 15 59561
rect -307 59240 -306 59560
rect 14 59240 15 59560
rect -307 59239 15 59240
rect -198 58841 -94 59239
rect 282 59188 302 59612
rect 366 59188 386 59612
rect 282 58892 386 59188
rect -307 58840 15 58841
rect -307 58520 -306 58840
rect 14 58520 15 58840
rect -307 58519 15 58520
rect -198 58121 -94 58519
rect 282 58468 302 58892
rect 366 58468 386 58892
rect 282 58172 386 58468
rect -307 58120 15 58121
rect -307 57800 -306 58120
rect 14 57800 15 58120
rect -307 57799 15 57800
rect -198 57401 -94 57799
rect 282 57748 302 58172
rect 366 57748 386 58172
rect 282 57452 386 57748
rect -307 57400 15 57401
rect -307 57080 -306 57400
rect 14 57080 15 57400
rect -307 57079 15 57080
rect -198 56681 -94 57079
rect 282 57028 302 57452
rect 366 57028 386 57452
rect 282 56732 386 57028
rect -307 56680 15 56681
rect -307 56360 -306 56680
rect 14 56360 15 56680
rect -307 56359 15 56360
rect -198 55961 -94 56359
rect 282 56308 302 56732
rect 366 56308 386 56732
rect 282 56012 386 56308
rect -307 55960 15 55961
rect -307 55640 -306 55960
rect 14 55640 15 55960
rect -307 55639 15 55640
rect -198 55241 -94 55639
rect 282 55588 302 56012
rect 366 55588 386 56012
rect 282 55292 386 55588
rect -307 55240 15 55241
rect -307 54920 -306 55240
rect 14 54920 15 55240
rect -307 54919 15 54920
rect -198 54521 -94 54919
rect 282 54868 302 55292
rect 366 54868 386 55292
rect 282 54572 386 54868
rect -307 54520 15 54521
rect -307 54200 -306 54520
rect 14 54200 15 54520
rect -307 54199 15 54200
rect -198 53801 -94 54199
rect 282 54148 302 54572
rect 366 54148 386 54572
rect 282 53852 386 54148
rect -307 53800 15 53801
rect -307 53480 -306 53800
rect 14 53480 15 53800
rect -307 53479 15 53480
rect -198 53081 -94 53479
rect 282 53428 302 53852
rect 366 53428 386 53852
rect 282 53132 386 53428
rect -307 53080 15 53081
rect -307 52760 -306 53080
rect 14 52760 15 53080
rect -307 52759 15 52760
rect -198 52361 -94 52759
rect 282 52708 302 53132
rect 366 52708 386 53132
rect 282 52412 386 52708
rect -307 52360 15 52361
rect -307 52040 -306 52360
rect 14 52040 15 52360
rect -307 52039 15 52040
rect -198 51641 -94 52039
rect 282 51988 302 52412
rect 366 51988 386 52412
rect 282 51692 386 51988
rect -307 51640 15 51641
rect -307 51320 -306 51640
rect 14 51320 15 51640
rect -307 51319 15 51320
rect -198 50921 -94 51319
rect 282 51268 302 51692
rect 366 51268 386 51692
rect 282 50972 386 51268
rect -307 50920 15 50921
rect -307 50600 -306 50920
rect 14 50600 15 50920
rect -307 50599 15 50600
rect -198 50201 -94 50599
rect 282 50548 302 50972
rect 366 50548 386 50972
rect 282 50252 386 50548
rect -307 50200 15 50201
rect -307 49880 -306 50200
rect 14 49880 15 50200
rect -307 49879 15 49880
rect -198 49481 -94 49879
rect 282 49828 302 50252
rect 366 49828 386 50252
rect 282 49532 386 49828
rect -307 49480 15 49481
rect -307 49160 -306 49480
rect 14 49160 15 49480
rect -307 49159 15 49160
rect -198 48761 -94 49159
rect 282 49108 302 49532
rect 366 49108 386 49532
rect 282 48812 386 49108
rect -307 48760 15 48761
rect -307 48440 -306 48760
rect 14 48440 15 48760
rect -307 48439 15 48440
rect -198 48041 -94 48439
rect 282 48388 302 48812
rect 366 48388 386 48812
rect 282 48092 386 48388
rect -307 48040 15 48041
rect -307 47720 -306 48040
rect 14 47720 15 48040
rect -307 47719 15 47720
rect -198 47321 -94 47719
rect 282 47668 302 48092
rect 366 47668 386 48092
rect 282 47372 386 47668
rect -307 47320 15 47321
rect -307 47000 -306 47320
rect 14 47000 15 47320
rect -307 46999 15 47000
rect -198 46601 -94 46999
rect 282 46948 302 47372
rect 366 46948 386 47372
rect 282 46652 386 46948
rect -307 46600 15 46601
rect -307 46280 -306 46600
rect 14 46280 15 46600
rect -307 46279 15 46280
rect -198 45881 -94 46279
rect 282 46228 302 46652
rect 366 46228 386 46652
rect 282 45932 386 46228
rect -307 45880 15 45881
rect -307 45560 -306 45880
rect 14 45560 15 45880
rect -307 45559 15 45560
rect -198 45161 -94 45559
rect 282 45508 302 45932
rect 366 45508 386 45932
rect 282 45212 386 45508
rect -307 45160 15 45161
rect -307 44840 -306 45160
rect 14 44840 15 45160
rect -307 44839 15 44840
rect -198 44441 -94 44839
rect 282 44788 302 45212
rect 366 44788 386 45212
rect 282 44492 386 44788
rect -307 44440 15 44441
rect -307 44120 -306 44440
rect 14 44120 15 44440
rect -307 44119 15 44120
rect -198 43721 -94 44119
rect 282 44068 302 44492
rect 366 44068 386 44492
rect 282 43772 386 44068
rect -307 43720 15 43721
rect -307 43400 -306 43720
rect 14 43400 15 43720
rect -307 43399 15 43400
rect -198 43001 -94 43399
rect 282 43348 302 43772
rect 366 43348 386 43772
rect 282 43052 386 43348
rect -307 43000 15 43001
rect -307 42680 -306 43000
rect 14 42680 15 43000
rect -307 42679 15 42680
rect -198 42281 -94 42679
rect 282 42628 302 43052
rect 366 42628 386 43052
rect 282 42332 386 42628
rect -307 42280 15 42281
rect -307 41960 -306 42280
rect 14 41960 15 42280
rect -307 41959 15 41960
rect -198 41561 -94 41959
rect 282 41908 302 42332
rect 366 41908 386 42332
rect 282 41612 386 41908
rect -307 41560 15 41561
rect -307 41240 -306 41560
rect 14 41240 15 41560
rect -307 41239 15 41240
rect -198 40841 -94 41239
rect 282 41188 302 41612
rect 366 41188 386 41612
rect 282 40892 386 41188
rect -307 40840 15 40841
rect -307 40520 -306 40840
rect 14 40520 15 40840
rect -307 40519 15 40520
rect -198 40121 -94 40519
rect 282 40468 302 40892
rect 366 40468 386 40892
rect 282 40172 386 40468
rect -307 40120 15 40121
rect -307 39800 -306 40120
rect 14 39800 15 40120
rect -307 39799 15 39800
rect -198 39401 -94 39799
rect 282 39748 302 40172
rect 366 39748 386 40172
rect 282 39452 386 39748
rect -307 39400 15 39401
rect -307 39080 -306 39400
rect 14 39080 15 39400
rect -307 39079 15 39080
rect -198 38681 -94 39079
rect 282 39028 302 39452
rect 366 39028 386 39452
rect 282 38732 386 39028
rect -307 38680 15 38681
rect -307 38360 -306 38680
rect 14 38360 15 38680
rect -307 38359 15 38360
rect -198 37961 -94 38359
rect 282 38308 302 38732
rect 366 38308 386 38732
rect 282 38012 386 38308
rect -307 37960 15 37961
rect -307 37640 -306 37960
rect 14 37640 15 37960
rect -307 37639 15 37640
rect -198 37241 -94 37639
rect 282 37588 302 38012
rect 366 37588 386 38012
rect 282 37292 386 37588
rect -307 37240 15 37241
rect -307 36920 -306 37240
rect 14 36920 15 37240
rect -307 36919 15 36920
rect -198 36521 -94 36919
rect 282 36868 302 37292
rect 366 36868 386 37292
rect 282 36572 386 36868
rect -307 36520 15 36521
rect -307 36200 -306 36520
rect 14 36200 15 36520
rect -307 36199 15 36200
rect -198 35801 -94 36199
rect 282 36148 302 36572
rect 366 36148 386 36572
rect 282 35852 386 36148
rect -307 35800 15 35801
rect -307 35480 -306 35800
rect 14 35480 15 35800
rect -307 35479 15 35480
rect -198 35081 -94 35479
rect 282 35428 302 35852
rect 366 35428 386 35852
rect 282 35132 386 35428
rect -307 35080 15 35081
rect -307 34760 -306 35080
rect 14 34760 15 35080
rect -307 34759 15 34760
rect -198 34361 -94 34759
rect 282 34708 302 35132
rect 366 34708 386 35132
rect 282 34412 386 34708
rect -307 34360 15 34361
rect -307 34040 -306 34360
rect 14 34040 15 34360
rect -307 34039 15 34040
rect -198 33641 -94 34039
rect 282 33988 302 34412
rect 366 33988 386 34412
rect 282 33692 386 33988
rect -307 33640 15 33641
rect -307 33320 -306 33640
rect 14 33320 15 33640
rect -307 33319 15 33320
rect -198 32921 -94 33319
rect 282 33268 302 33692
rect 366 33268 386 33692
rect 282 32972 386 33268
rect -307 32920 15 32921
rect -307 32600 -306 32920
rect 14 32600 15 32920
rect -307 32599 15 32600
rect -198 32201 -94 32599
rect 282 32548 302 32972
rect 366 32548 386 32972
rect 282 32252 386 32548
rect -307 32200 15 32201
rect -307 31880 -306 32200
rect 14 31880 15 32200
rect -307 31879 15 31880
rect -198 31481 -94 31879
rect 282 31828 302 32252
rect 366 31828 386 32252
rect 282 31532 386 31828
rect -307 31480 15 31481
rect -307 31160 -306 31480
rect 14 31160 15 31480
rect -307 31159 15 31160
rect -198 30761 -94 31159
rect 282 31108 302 31532
rect 366 31108 386 31532
rect 282 30812 386 31108
rect -307 30760 15 30761
rect -307 30440 -306 30760
rect 14 30440 15 30760
rect -307 30439 15 30440
rect -198 30041 -94 30439
rect 282 30388 302 30812
rect 366 30388 386 30812
rect 282 30092 386 30388
rect -307 30040 15 30041
rect -307 29720 -306 30040
rect 14 29720 15 30040
rect -307 29719 15 29720
rect -198 29321 -94 29719
rect 282 29668 302 30092
rect 366 29668 386 30092
rect 282 29372 386 29668
rect -307 29320 15 29321
rect -307 29000 -306 29320
rect 14 29000 15 29320
rect -307 28999 15 29000
rect -198 28601 -94 28999
rect 282 28948 302 29372
rect 366 28948 386 29372
rect 282 28652 386 28948
rect -307 28600 15 28601
rect -307 28280 -306 28600
rect 14 28280 15 28600
rect -307 28279 15 28280
rect -198 27881 -94 28279
rect 282 28228 302 28652
rect 366 28228 386 28652
rect 282 27932 386 28228
rect -307 27880 15 27881
rect -307 27560 -306 27880
rect 14 27560 15 27880
rect -307 27559 15 27560
rect -198 27161 -94 27559
rect 282 27508 302 27932
rect 366 27508 386 27932
rect 282 27212 386 27508
rect -307 27160 15 27161
rect -307 26840 -306 27160
rect 14 26840 15 27160
rect -307 26839 15 26840
rect -198 26441 -94 26839
rect 282 26788 302 27212
rect 366 26788 386 27212
rect 282 26492 386 26788
rect -307 26440 15 26441
rect -307 26120 -306 26440
rect 14 26120 15 26440
rect -307 26119 15 26120
rect -198 25721 -94 26119
rect 282 26068 302 26492
rect 366 26068 386 26492
rect 282 25772 386 26068
rect -307 25720 15 25721
rect -307 25400 -306 25720
rect 14 25400 15 25720
rect -307 25399 15 25400
rect -198 25001 -94 25399
rect 282 25348 302 25772
rect 366 25348 386 25772
rect 282 25052 386 25348
rect -307 25000 15 25001
rect -307 24680 -306 25000
rect 14 24680 15 25000
rect -307 24679 15 24680
rect -198 24281 -94 24679
rect 282 24628 302 25052
rect 366 24628 386 25052
rect 282 24332 386 24628
rect -307 24280 15 24281
rect -307 23960 -306 24280
rect 14 23960 15 24280
rect -307 23959 15 23960
rect -198 23561 -94 23959
rect 282 23908 302 24332
rect 366 23908 386 24332
rect 282 23612 386 23908
rect -307 23560 15 23561
rect -307 23240 -306 23560
rect 14 23240 15 23560
rect -307 23239 15 23240
rect -198 22841 -94 23239
rect 282 23188 302 23612
rect 366 23188 386 23612
rect 282 22892 386 23188
rect -307 22840 15 22841
rect -307 22520 -306 22840
rect 14 22520 15 22840
rect -307 22519 15 22520
rect -198 22121 -94 22519
rect 282 22468 302 22892
rect 366 22468 386 22892
rect 282 22172 386 22468
rect -307 22120 15 22121
rect -307 21800 -306 22120
rect 14 21800 15 22120
rect -307 21799 15 21800
rect -198 21401 -94 21799
rect 282 21748 302 22172
rect 366 21748 386 22172
rect 282 21452 386 21748
rect -307 21400 15 21401
rect -307 21080 -306 21400
rect 14 21080 15 21400
rect -307 21079 15 21080
rect -198 20681 -94 21079
rect 282 21028 302 21452
rect 366 21028 386 21452
rect 282 20732 386 21028
rect -307 20680 15 20681
rect -307 20360 -306 20680
rect 14 20360 15 20680
rect -307 20359 15 20360
rect -198 19961 -94 20359
rect 282 20308 302 20732
rect 366 20308 386 20732
rect 282 20012 386 20308
rect -307 19960 15 19961
rect -307 19640 -306 19960
rect 14 19640 15 19960
rect -307 19639 15 19640
rect -198 19241 -94 19639
rect 282 19588 302 20012
rect 366 19588 386 20012
rect 282 19292 386 19588
rect -307 19240 15 19241
rect -307 18920 -306 19240
rect 14 18920 15 19240
rect -307 18919 15 18920
rect -198 18521 -94 18919
rect 282 18868 302 19292
rect 366 18868 386 19292
rect 282 18572 386 18868
rect -307 18520 15 18521
rect -307 18200 -306 18520
rect 14 18200 15 18520
rect -307 18199 15 18200
rect -198 17801 -94 18199
rect 282 18148 302 18572
rect 366 18148 386 18572
rect 282 17852 386 18148
rect -307 17800 15 17801
rect -307 17480 -306 17800
rect 14 17480 15 17800
rect -307 17479 15 17480
rect -198 17081 -94 17479
rect 282 17428 302 17852
rect 366 17428 386 17852
rect 282 17132 386 17428
rect -307 17080 15 17081
rect -307 16760 -306 17080
rect 14 16760 15 17080
rect -307 16759 15 16760
rect -198 16361 -94 16759
rect 282 16708 302 17132
rect 366 16708 386 17132
rect 282 16412 386 16708
rect -307 16360 15 16361
rect -307 16040 -306 16360
rect 14 16040 15 16360
rect -307 16039 15 16040
rect -198 15641 -94 16039
rect 282 15988 302 16412
rect 366 15988 386 16412
rect 282 15692 386 15988
rect -307 15640 15 15641
rect -307 15320 -306 15640
rect 14 15320 15 15640
rect -307 15319 15 15320
rect -198 14921 -94 15319
rect 282 15268 302 15692
rect 366 15268 386 15692
rect 282 14972 386 15268
rect -307 14920 15 14921
rect -307 14600 -306 14920
rect 14 14600 15 14920
rect -307 14599 15 14600
rect -198 14201 -94 14599
rect 282 14548 302 14972
rect 366 14548 386 14972
rect 282 14252 386 14548
rect -307 14200 15 14201
rect -307 13880 -306 14200
rect 14 13880 15 14200
rect -307 13879 15 13880
rect -198 13481 -94 13879
rect 282 13828 302 14252
rect 366 13828 386 14252
rect 282 13532 386 13828
rect -307 13480 15 13481
rect -307 13160 -306 13480
rect 14 13160 15 13480
rect -307 13159 15 13160
rect -198 12761 -94 13159
rect 282 13108 302 13532
rect 366 13108 386 13532
rect 282 12812 386 13108
rect -307 12760 15 12761
rect -307 12440 -306 12760
rect 14 12440 15 12760
rect -307 12439 15 12440
rect -198 12041 -94 12439
rect 282 12388 302 12812
rect 366 12388 386 12812
rect 282 12092 386 12388
rect -307 12040 15 12041
rect -307 11720 -306 12040
rect 14 11720 15 12040
rect -307 11719 15 11720
rect -198 11321 -94 11719
rect 282 11668 302 12092
rect 366 11668 386 12092
rect 282 11372 386 11668
rect -307 11320 15 11321
rect -307 11000 -306 11320
rect 14 11000 15 11320
rect -307 10999 15 11000
rect -198 10601 -94 10999
rect 282 10948 302 11372
rect 366 10948 386 11372
rect 282 10652 386 10948
rect -307 10600 15 10601
rect -307 10280 -306 10600
rect 14 10280 15 10600
rect -307 10279 15 10280
rect -198 9881 -94 10279
rect 282 10228 302 10652
rect 366 10228 386 10652
rect 282 9932 386 10228
rect -307 9880 15 9881
rect -307 9560 -306 9880
rect 14 9560 15 9880
rect -307 9559 15 9560
rect -198 9161 -94 9559
rect 282 9508 302 9932
rect 366 9508 386 9932
rect 282 9212 386 9508
rect -307 9160 15 9161
rect -307 8840 -306 9160
rect 14 8840 15 9160
rect -307 8839 15 8840
rect -198 8441 -94 8839
rect 282 8788 302 9212
rect 366 8788 386 9212
rect 282 8492 386 8788
rect -307 8440 15 8441
rect -307 8120 -306 8440
rect 14 8120 15 8440
rect -307 8119 15 8120
rect -198 7721 -94 8119
rect 282 8068 302 8492
rect 366 8068 386 8492
rect 282 7772 386 8068
rect -307 7720 15 7721
rect -307 7400 -306 7720
rect 14 7400 15 7720
rect -307 7399 15 7400
rect -198 7001 -94 7399
rect 282 7348 302 7772
rect 366 7348 386 7772
rect 282 7052 386 7348
rect -307 7000 15 7001
rect -307 6680 -306 7000
rect 14 6680 15 7000
rect -307 6679 15 6680
rect -198 6281 -94 6679
rect 282 6628 302 7052
rect 366 6628 386 7052
rect 282 6332 386 6628
rect -307 6280 15 6281
rect -307 5960 -306 6280
rect 14 5960 15 6280
rect -307 5959 15 5960
rect -198 5561 -94 5959
rect 282 5908 302 6332
rect 366 5908 386 6332
rect 282 5612 386 5908
rect -307 5560 15 5561
rect -307 5240 -306 5560
rect 14 5240 15 5560
rect -307 5239 15 5240
rect -198 4841 -94 5239
rect 282 5188 302 5612
rect 366 5188 386 5612
rect 282 4892 386 5188
rect -307 4840 15 4841
rect -307 4520 -306 4840
rect 14 4520 15 4840
rect -307 4519 15 4520
rect -198 4121 -94 4519
rect 282 4468 302 4892
rect 366 4468 386 4892
rect 282 4172 386 4468
rect -307 4120 15 4121
rect -307 3800 -306 4120
rect 14 3800 15 4120
rect -307 3799 15 3800
rect -198 3401 -94 3799
rect 282 3748 302 4172
rect 366 3748 386 4172
rect 282 3452 386 3748
rect -307 3400 15 3401
rect -307 3080 -306 3400
rect 14 3080 15 3400
rect -307 3079 15 3080
rect -198 2681 -94 3079
rect 282 3028 302 3452
rect 366 3028 386 3452
rect 282 2732 386 3028
rect -307 2680 15 2681
rect -307 2360 -306 2680
rect 14 2360 15 2680
rect -307 2359 15 2360
rect -198 1961 -94 2359
rect 282 2308 302 2732
rect 366 2308 386 2732
rect 282 2012 386 2308
rect -307 1960 15 1961
rect -307 1640 -306 1960
rect 14 1640 15 1960
rect -307 1639 15 1640
rect -198 1241 -94 1639
rect 282 1588 302 2012
rect 366 1588 386 2012
rect 282 1292 386 1588
rect -307 1240 15 1241
rect -307 920 -306 1240
rect 14 920 15 1240
rect -307 919 15 920
rect -198 521 -94 919
rect 282 868 302 1292
rect 366 868 386 1292
rect 282 572 386 868
rect -307 520 15 521
rect -307 200 -306 520
rect 14 200 15 520
rect -307 199 15 200
rect -198 -199 -94 199
rect 282 148 302 572
rect 366 148 386 572
rect 282 -148 386 148
rect -307 -200 15 -199
rect -307 -520 -306 -200
rect 14 -520 15 -200
rect -307 -521 15 -520
rect -198 -919 -94 -521
rect 282 -572 302 -148
rect 366 -572 386 -148
rect 282 -868 386 -572
rect -307 -920 15 -919
rect -307 -1240 -306 -920
rect 14 -1240 15 -920
rect -307 -1241 15 -1240
rect -198 -1639 -94 -1241
rect 282 -1292 302 -868
rect 366 -1292 386 -868
rect 282 -1588 386 -1292
rect -307 -1640 15 -1639
rect -307 -1960 -306 -1640
rect 14 -1960 15 -1640
rect -307 -1961 15 -1960
rect -198 -2359 -94 -1961
rect 282 -2012 302 -1588
rect 366 -2012 386 -1588
rect 282 -2308 386 -2012
rect -307 -2360 15 -2359
rect -307 -2680 -306 -2360
rect 14 -2680 15 -2360
rect -307 -2681 15 -2680
rect -198 -3079 -94 -2681
rect 282 -2732 302 -2308
rect 366 -2732 386 -2308
rect 282 -3028 386 -2732
rect -307 -3080 15 -3079
rect -307 -3400 -306 -3080
rect 14 -3400 15 -3080
rect -307 -3401 15 -3400
rect -198 -3799 -94 -3401
rect 282 -3452 302 -3028
rect 366 -3452 386 -3028
rect 282 -3748 386 -3452
rect -307 -3800 15 -3799
rect -307 -4120 -306 -3800
rect 14 -4120 15 -3800
rect -307 -4121 15 -4120
rect -198 -4519 -94 -4121
rect 282 -4172 302 -3748
rect 366 -4172 386 -3748
rect 282 -4468 386 -4172
rect -307 -4520 15 -4519
rect -307 -4840 -306 -4520
rect 14 -4840 15 -4520
rect -307 -4841 15 -4840
rect -198 -5239 -94 -4841
rect 282 -4892 302 -4468
rect 366 -4892 386 -4468
rect 282 -5188 386 -4892
rect -307 -5240 15 -5239
rect -307 -5560 -306 -5240
rect 14 -5560 15 -5240
rect -307 -5561 15 -5560
rect -198 -5959 -94 -5561
rect 282 -5612 302 -5188
rect 366 -5612 386 -5188
rect 282 -5908 386 -5612
rect -307 -5960 15 -5959
rect -307 -6280 -306 -5960
rect 14 -6280 15 -5960
rect -307 -6281 15 -6280
rect -198 -6679 -94 -6281
rect 282 -6332 302 -5908
rect 366 -6332 386 -5908
rect 282 -6628 386 -6332
rect -307 -6680 15 -6679
rect -307 -7000 -306 -6680
rect 14 -7000 15 -6680
rect -307 -7001 15 -7000
rect -198 -7399 -94 -7001
rect 282 -7052 302 -6628
rect 366 -7052 386 -6628
rect 282 -7348 386 -7052
rect -307 -7400 15 -7399
rect -307 -7720 -306 -7400
rect 14 -7720 15 -7400
rect -307 -7721 15 -7720
rect -198 -8119 -94 -7721
rect 282 -7772 302 -7348
rect 366 -7772 386 -7348
rect 282 -8068 386 -7772
rect -307 -8120 15 -8119
rect -307 -8440 -306 -8120
rect 14 -8440 15 -8120
rect -307 -8441 15 -8440
rect -198 -8839 -94 -8441
rect 282 -8492 302 -8068
rect 366 -8492 386 -8068
rect 282 -8788 386 -8492
rect -307 -8840 15 -8839
rect -307 -9160 -306 -8840
rect 14 -9160 15 -8840
rect -307 -9161 15 -9160
rect -198 -9559 -94 -9161
rect 282 -9212 302 -8788
rect 366 -9212 386 -8788
rect 282 -9508 386 -9212
rect -307 -9560 15 -9559
rect -307 -9880 -306 -9560
rect 14 -9880 15 -9560
rect -307 -9881 15 -9880
rect -198 -10279 -94 -9881
rect 282 -9932 302 -9508
rect 366 -9932 386 -9508
rect 282 -10228 386 -9932
rect -307 -10280 15 -10279
rect -307 -10600 -306 -10280
rect 14 -10600 15 -10280
rect -307 -10601 15 -10600
rect -198 -10999 -94 -10601
rect 282 -10652 302 -10228
rect 366 -10652 386 -10228
rect 282 -10948 386 -10652
rect -307 -11000 15 -10999
rect -307 -11320 -306 -11000
rect 14 -11320 15 -11000
rect -307 -11321 15 -11320
rect -198 -11719 -94 -11321
rect 282 -11372 302 -10948
rect 366 -11372 386 -10948
rect 282 -11668 386 -11372
rect -307 -11720 15 -11719
rect -307 -12040 -306 -11720
rect 14 -12040 15 -11720
rect -307 -12041 15 -12040
rect -198 -12439 -94 -12041
rect 282 -12092 302 -11668
rect 366 -12092 386 -11668
rect 282 -12388 386 -12092
rect -307 -12440 15 -12439
rect -307 -12760 -306 -12440
rect 14 -12760 15 -12440
rect -307 -12761 15 -12760
rect -198 -13159 -94 -12761
rect 282 -12812 302 -12388
rect 366 -12812 386 -12388
rect 282 -13108 386 -12812
rect -307 -13160 15 -13159
rect -307 -13480 -306 -13160
rect 14 -13480 15 -13160
rect -307 -13481 15 -13480
rect -198 -13879 -94 -13481
rect 282 -13532 302 -13108
rect 366 -13532 386 -13108
rect 282 -13828 386 -13532
rect -307 -13880 15 -13879
rect -307 -14200 -306 -13880
rect 14 -14200 15 -13880
rect -307 -14201 15 -14200
rect -198 -14599 -94 -14201
rect 282 -14252 302 -13828
rect 366 -14252 386 -13828
rect 282 -14548 386 -14252
rect -307 -14600 15 -14599
rect -307 -14920 -306 -14600
rect 14 -14920 15 -14600
rect -307 -14921 15 -14920
rect -198 -15319 -94 -14921
rect 282 -14972 302 -14548
rect 366 -14972 386 -14548
rect 282 -15268 386 -14972
rect -307 -15320 15 -15319
rect -307 -15640 -306 -15320
rect 14 -15640 15 -15320
rect -307 -15641 15 -15640
rect -198 -16039 -94 -15641
rect 282 -15692 302 -15268
rect 366 -15692 386 -15268
rect 282 -15988 386 -15692
rect -307 -16040 15 -16039
rect -307 -16360 -306 -16040
rect 14 -16360 15 -16040
rect -307 -16361 15 -16360
rect -198 -16759 -94 -16361
rect 282 -16412 302 -15988
rect 366 -16412 386 -15988
rect 282 -16708 386 -16412
rect -307 -16760 15 -16759
rect -307 -17080 -306 -16760
rect 14 -17080 15 -16760
rect -307 -17081 15 -17080
rect -198 -17479 -94 -17081
rect 282 -17132 302 -16708
rect 366 -17132 386 -16708
rect 282 -17428 386 -17132
rect -307 -17480 15 -17479
rect -307 -17800 -306 -17480
rect 14 -17800 15 -17480
rect -307 -17801 15 -17800
rect -198 -18199 -94 -17801
rect 282 -17852 302 -17428
rect 366 -17852 386 -17428
rect 282 -18148 386 -17852
rect -307 -18200 15 -18199
rect -307 -18520 -306 -18200
rect 14 -18520 15 -18200
rect -307 -18521 15 -18520
rect -198 -18919 -94 -18521
rect 282 -18572 302 -18148
rect 366 -18572 386 -18148
rect 282 -18868 386 -18572
rect -307 -18920 15 -18919
rect -307 -19240 -306 -18920
rect 14 -19240 15 -18920
rect -307 -19241 15 -19240
rect -198 -19639 -94 -19241
rect 282 -19292 302 -18868
rect 366 -19292 386 -18868
rect 282 -19588 386 -19292
rect -307 -19640 15 -19639
rect -307 -19960 -306 -19640
rect 14 -19960 15 -19640
rect -307 -19961 15 -19960
rect -198 -20359 -94 -19961
rect 282 -20012 302 -19588
rect 366 -20012 386 -19588
rect 282 -20308 386 -20012
rect -307 -20360 15 -20359
rect -307 -20680 -306 -20360
rect 14 -20680 15 -20360
rect -307 -20681 15 -20680
rect -198 -21079 -94 -20681
rect 282 -20732 302 -20308
rect 366 -20732 386 -20308
rect 282 -21028 386 -20732
rect -307 -21080 15 -21079
rect -307 -21400 -306 -21080
rect 14 -21400 15 -21080
rect -307 -21401 15 -21400
rect -198 -21799 -94 -21401
rect 282 -21452 302 -21028
rect 366 -21452 386 -21028
rect 282 -21748 386 -21452
rect -307 -21800 15 -21799
rect -307 -22120 -306 -21800
rect 14 -22120 15 -21800
rect -307 -22121 15 -22120
rect -198 -22519 -94 -22121
rect 282 -22172 302 -21748
rect 366 -22172 386 -21748
rect 282 -22468 386 -22172
rect -307 -22520 15 -22519
rect -307 -22840 -306 -22520
rect 14 -22840 15 -22520
rect -307 -22841 15 -22840
rect -198 -23239 -94 -22841
rect 282 -22892 302 -22468
rect 366 -22892 386 -22468
rect 282 -23188 386 -22892
rect -307 -23240 15 -23239
rect -307 -23560 -306 -23240
rect 14 -23560 15 -23240
rect -307 -23561 15 -23560
rect -198 -23959 -94 -23561
rect 282 -23612 302 -23188
rect 366 -23612 386 -23188
rect 282 -23908 386 -23612
rect -307 -23960 15 -23959
rect -307 -24280 -306 -23960
rect 14 -24280 15 -23960
rect -307 -24281 15 -24280
rect -198 -24679 -94 -24281
rect 282 -24332 302 -23908
rect 366 -24332 386 -23908
rect 282 -24628 386 -24332
rect -307 -24680 15 -24679
rect -307 -25000 -306 -24680
rect 14 -25000 15 -24680
rect -307 -25001 15 -25000
rect -198 -25399 -94 -25001
rect 282 -25052 302 -24628
rect 366 -25052 386 -24628
rect 282 -25348 386 -25052
rect -307 -25400 15 -25399
rect -307 -25720 -306 -25400
rect 14 -25720 15 -25400
rect -307 -25721 15 -25720
rect -198 -26119 -94 -25721
rect 282 -25772 302 -25348
rect 366 -25772 386 -25348
rect 282 -26068 386 -25772
rect -307 -26120 15 -26119
rect -307 -26440 -306 -26120
rect 14 -26440 15 -26120
rect -307 -26441 15 -26440
rect -198 -26839 -94 -26441
rect 282 -26492 302 -26068
rect 366 -26492 386 -26068
rect 282 -26788 386 -26492
rect -307 -26840 15 -26839
rect -307 -27160 -306 -26840
rect 14 -27160 15 -26840
rect -307 -27161 15 -27160
rect -198 -27559 -94 -27161
rect 282 -27212 302 -26788
rect 366 -27212 386 -26788
rect 282 -27508 386 -27212
rect -307 -27560 15 -27559
rect -307 -27880 -306 -27560
rect 14 -27880 15 -27560
rect -307 -27881 15 -27880
rect -198 -28279 -94 -27881
rect 282 -27932 302 -27508
rect 366 -27932 386 -27508
rect 282 -28228 386 -27932
rect -307 -28280 15 -28279
rect -307 -28600 -306 -28280
rect 14 -28600 15 -28280
rect -307 -28601 15 -28600
rect -198 -28999 -94 -28601
rect 282 -28652 302 -28228
rect 366 -28652 386 -28228
rect 282 -28948 386 -28652
rect -307 -29000 15 -28999
rect -307 -29320 -306 -29000
rect 14 -29320 15 -29000
rect -307 -29321 15 -29320
rect -198 -29719 -94 -29321
rect 282 -29372 302 -28948
rect 366 -29372 386 -28948
rect 282 -29668 386 -29372
rect -307 -29720 15 -29719
rect -307 -30040 -306 -29720
rect 14 -30040 15 -29720
rect -307 -30041 15 -30040
rect -198 -30439 -94 -30041
rect 282 -30092 302 -29668
rect 366 -30092 386 -29668
rect 282 -30388 386 -30092
rect -307 -30440 15 -30439
rect -307 -30760 -306 -30440
rect 14 -30760 15 -30440
rect -307 -30761 15 -30760
rect -198 -31159 -94 -30761
rect 282 -30812 302 -30388
rect 366 -30812 386 -30388
rect 282 -31108 386 -30812
rect -307 -31160 15 -31159
rect -307 -31480 -306 -31160
rect 14 -31480 15 -31160
rect -307 -31481 15 -31480
rect -198 -31879 -94 -31481
rect 282 -31532 302 -31108
rect 366 -31532 386 -31108
rect 282 -31828 386 -31532
rect -307 -31880 15 -31879
rect -307 -32200 -306 -31880
rect 14 -32200 15 -31880
rect -307 -32201 15 -32200
rect -198 -32599 -94 -32201
rect 282 -32252 302 -31828
rect 366 -32252 386 -31828
rect 282 -32548 386 -32252
rect -307 -32600 15 -32599
rect -307 -32920 -306 -32600
rect 14 -32920 15 -32600
rect -307 -32921 15 -32920
rect -198 -33319 -94 -32921
rect 282 -32972 302 -32548
rect 366 -32972 386 -32548
rect 282 -33268 386 -32972
rect -307 -33320 15 -33319
rect -307 -33640 -306 -33320
rect 14 -33640 15 -33320
rect -307 -33641 15 -33640
rect -198 -34039 -94 -33641
rect 282 -33692 302 -33268
rect 366 -33692 386 -33268
rect 282 -33988 386 -33692
rect -307 -34040 15 -34039
rect -307 -34360 -306 -34040
rect 14 -34360 15 -34040
rect -307 -34361 15 -34360
rect -198 -34759 -94 -34361
rect 282 -34412 302 -33988
rect 366 -34412 386 -33988
rect 282 -34708 386 -34412
rect -307 -34760 15 -34759
rect -307 -35080 -306 -34760
rect 14 -35080 15 -34760
rect -307 -35081 15 -35080
rect -198 -35479 -94 -35081
rect 282 -35132 302 -34708
rect 366 -35132 386 -34708
rect 282 -35428 386 -35132
rect -307 -35480 15 -35479
rect -307 -35800 -306 -35480
rect 14 -35800 15 -35480
rect -307 -35801 15 -35800
rect -198 -36199 -94 -35801
rect 282 -35852 302 -35428
rect 366 -35852 386 -35428
rect 282 -36148 386 -35852
rect -307 -36200 15 -36199
rect -307 -36520 -306 -36200
rect 14 -36520 15 -36200
rect -307 -36521 15 -36520
rect -198 -36919 -94 -36521
rect 282 -36572 302 -36148
rect 366 -36572 386 -36148
rect 282 -36868 386 -36572
rect -307 -36920 15 -36919
rect -307 -37240 -306 -36920
rect 14 -37240 15 -36920
rect -307 -37241 15 -37240
rect -198 -37639 -94 -37241
rect 282 -37292 302 -36868
rect 366 -37292 386 -36868
rect 282 -37588 386 -37292
rect -307 -37640 15 -37639
rect -307 -37960 -306 -37640
rect 14 -37960 15 -37640
rect -307 -37961 15 -37960
rect -198 -38359 -94 -37961
rect 282 -38012 302 -37588
rect 366 -38012 386 -37588
rect 282 -38308 386 -38012
rect -307 -38360 15 -38359
rect -307 -38680 -306 -38360
rect 14 -38680 15 -38360
rect -307 -38681 15 -38680
rect -198 -39079 -94 -38681
rect 282 -38732 302 -38308
rect 366 -38732 386 -38308
rect 282 -39028 386 -38732
rect -307 -39080 15 -39079
rect -307 -39400 -306 -39080
rect 14 -39400 15 -39080
rect -307 -39401 15 -39400
rect -198 -39799 -94 -39401
rect 282 -39452 302 -39028
rect 366 -39452 386 -39028
rect 282 -39748 386 -39452
rect -307 -39800 15 -39799
rect -307 -40120 -306 -39800
rect 14 -40120 15 -39800
rect -307 -40121 15 -40120
rect -198 -40519 -94 -40121
rect 282 -40172 302 -39748
rect 366 -40172 386 -39748
rect 282 -40468 386 -40172
rect -307 -40520 15 -40519
rect -307 -40840 -306 -40520
rect 14 -40840 15 -40520
rect -307 -40841 15 -40840
rect -198 -41239 -94 -40841
rect 282 -40892 302 -40468
rect 366 -40892 386 -40468
rect 282 -41188 386 -40892
rect -307 -41240 15 -41239
rect -307 -41560 -306 -41240
rect 14 -41560 15 -41240
rect -307 -41561 15 -41560
rect -198 -41959 -94 -41561
rect 282 -41612 302 -41188
rect 366 -41612 386 -41188
rect 282 -41908 386 -41612
rect -307 -41960 15 -41959
rect -307 -42280 -306 -41960
rect 14 -42280 15 -41960
rect -307 -42281 15 -42280
rect -198 -42679 -94 -42281
rect 282 -42332 302 -41908
rect 366 -42332 386 -41908
rect 282 -42628 386 -42332
rect -307 -42680 15 -42679
rect -307 -43000 -306 -42680
rect 14 -43000 15 -42680
rect -307 -43001 15 -43000
rect -198 -43399 -94 -43001
rect 282 -43052 302 -42628
rect 366 -43052 386 -42628
rect 282 -43348 386 -43052
rect -307 -43400 15 -43399
rect -307 -43720 -306 -43400
rect 14 -43720 15 -43400
rect -307 -43721 15 -43720
rect -198 -44119 -94 -43721
rect 282 -43772 302 -43348
rect 366 -43772 386 -43348
rect 282 -44068 386 -43772
rect -307 -44120 15 -44119
rect -307 -44440 -306 -44120
rect 14 -44440 15 -44120
rect -307 -44441 15 -44440
rect -198 -44839 -94 -44441
rect 282 -44492 302 -44068
rect 366 -44492 386 -44068
rect 282 -44788 386 -44492
rect -307 -44840 15 -44839
rect -307 -45160 -306 -44840
rect 14 -45160 15 -44840
rect -307 -45161 15 -45160
rect -198 -45559 -94 -45161
rect 282 -45212 302 -44788
rect 366 -45212 386 -44788
rect 282 -45508 386 -45212
rect -307 -45560 15 -45559
rect -307 -45880 -306 -45560
rect 14 -45880 15 -45560
rect -307 -45881 15 -45880
rect -198 -46279 -94 -45881
rect 282 -45932 302 -45508
rect 366 -45932 386 -45508
rect 282 -46228 386 -45932
rect -307 -46280 15 -46279
rect -307 -46600 -306 -46280
rect 14 -46600 15 -46280
rect -307 -46601 15 -46600
rect -198 -46999 -94 -46601
rect 282 -46652 302 -46228
rect 366 -46652 386 -46228
rect 282 -46948 386 -46652
rect -307 -47000 15 -46999
rect -307 -47320 -306 -47000
rect 14 -47320 15 -47000
rect -307 -47321 15 -47320
rect -198 -47719 -94 -47321
rect 282 -47372 302 -46948
rect 366 -47372 386 -46948
rect 282 -47668 386 -47372
rect -307 -47720 15 -47719
rect -307 -48040 -306 -47720
rect 14 -48040 15 -47720
rect -307 -48041 15 -48040
rect -198 -48439 -94 -48041
rect 282 -48092 302 -47668
rect 366 -48092 386 -47668
rect 282 -48388 386 -48092
rect -307 -48440 15 -48439
rect -307 -48760 -306 -48440
rect 14 -48760 15 -48440
rect -307 -48761 15 -48760
rect -198 -49159 -94 -48761
rect 282 -48812 302 -48388
rect 366 -48812 386 -48388
rect 282 -49108 386 -48812
rect -307 -49160 15 -49159
rect -307 -49480 -306 -49160
rect 14 -49480 15 -49160
rect -307 -49481 15 -49480
rect -198 -49879 -94 -49481
rect 282 -49532 302 -49108
rect 366 -49532 386 -49108
rect 282 -49828 386 -49532
rect -307 -49880 15 -49879
rect -307 -50200 -306 -49880
rect 14 -50200 15 -49880
rect -307 -50201 15 -50200
rect -198 -50599 -94 -50201
rect 282 -50252 302 -49828
rect 366 -50252 386 -49828
rect 282 -50548 386 -50252
rect -307 -50600 15 -50599
rect -307 -50920 -306 -50600
rect 14 -50920 15 -50600
rect -307 -50921 15 -50920
rect -198 -51319 -94 -50921
rect 282 -50972 302 -50548
rect 366 -50972 386 -50548
rect 282 -51268 386 -50972
rect -307 -51320 15 -51319
rect -307 -51640 -306 -51320
rect 14 -51640 15 -51320
rect -307 -51641 15 -51640
rect -198 -52039 -94 -51641
rect 282 -51692 302 -51268
rect 366 -51692 386 -51268
rect 282 -51988 386 -51692
rect -307 -52040 15 -52039
rect -307 -52360 -306 -52040
rect 14 -52360 15 -52040
rect -307 -52361 15 -52360
rect -198 -52759 -94 -52361
rect 282 -52412 302 -51988
rect 366 -52412 386 -51988
rect 282 -52708 386 -52412
rect -307 -52760 15 -52759
rect -307 -53080 -306 -52760
rect 14 -53080 15 -52760
rect -307 -53081 15 -53080
rect -198 -53479 -94 -53081
rect 282 -53132 302 -52708
rect 366 -53132 386 -52708
rect 282 -53428 386 -53132
rect -307 -53480 15 -53479
rect -307 -53800 -306 -53480
rect 14 -53800 15 -53480
rect -307 -53801 15 -53800
rect -198 -54199 -94 -53801
rect 282 -53852 302 -53428
rect 366 -53852 386 -53428
rect 282 -54148 386 -53852
rect -307 -54200 15 -54199
rect -307 -54520 -306 -54200
rect 14 -54520 15 -54200
rect -307 -54521 15 -54520
rect -198 -54919 -94 -54521
rect 282 -54572 302 -54148
rect 366 -54572 386 -54148
rect 282 -54868 386 -54572
rect -307 -54920 15 -54919
rect -307 -55240 -306 -54920
rect 14 -55240 15 -54920
rect -307 -55241 15 -55240
rect -198 -55639 -94 -55241
rect 282 -55292 302 -54868
rect 366 -55292 386 -54868
rect 282 -55588 386 -55292
rect -307 -55640 15 -55639
rect -307 -55960 -306 -55640
rect 14 -55960 15 -55640
rect -307 -55961 15 -55960
rect -198 -56359 -94 -55961
rect 282 -56012 302 -55588
rect 366 -56012 386 -55588
rect 282 -56308 386 -56012
rect -307 -56360 15 -56359
rect -307 -56680 -306 -56360
rect 14 -56680 15 -56360
rect -307 -56681 15 -56680
rect -198 -57079 -94 -56681
rect 282 -56732 302 -56308
rect 366 -56732 386 -56308
rect 282 -57028 386 -56732
rect -307 -57080 15 -57079
rect -307 -57400 -306 -57080
rect 14 -57400 15 -57080
rect -307 -57401 15 -57400
rect -198 -57799 -94 -57401
rect 282 -57452 302 -57028
rect 366 -57452 386 -57028
rect 282 -57748 386 -57452
rect -307 -57800 15 -57799
rect -307 -58120 -306 -57800
rect 14 -58120 15 -57800
rect -307 -58121 15 -58120
rect -198 -58519 -94 -58121
rect 282 -58172 302 -57748
rect 366 -58172 386 -57748
rect 282 -58468 386 -58172
rect -307 -58520 15 -58519
rect -307 -58840 -306 -58520
rect 14 -58840 15 -58520
rect -307 -58841 15 -58840
rect -198 -59239 -94 -58841
rect 282 -58892 302 -58468
rect 366 -58892 386 -58468
rect 282 -59188 386 -58892
rect -307 -59240 15 -59239
rect -307 -59560 -306 -59240
rect 14 -59560 15 -59240
rect -307 -59561 15 -59560
rect -198 -59959 -94 -59561
rect 282 -59612 302 -59188
rect 366 -59612 386 -59188
rect 282 -59908 386 -59612
rect -307 -59960 15 -59959
rect -307 -60280 -306 -59960
rect 14 -60280 15 -59960
rect -307 -60281 15 -60280
rect -198 -60679 -94 -60281
rect 282 -60332 302 -59908
rect 366 -60332 386 -59908
rect 282 -60628 386 -60332
rect -307 -60680 15 -60679
rect -307 -61000 -306 -60680
rect 14 -61000 15 -60680
rect -307 -61001 15 -61000
rect -198 -61399 -94 -61001
rect 282 -61052 302 -60628
rect 366 -61052 386 -60628
rect 282 -61348 386 -61052
rect -307 -61400 15 -61399
rect -307 -61720 -306 -61400
rect 14 -61720 15 -61400
rect -307 -61721 15 -61720
rect -198 -62119 -94 -61721
rect 282 -61772 302 -61348
rect 366 -61772 386 -61348
rect 282 -62068 386 -61772
rect -307 -62120 15 -62119
rect -307 -62440 -306 -62120
rect 14 -62440 15 -62120
rect -307 -62441 15 -62440
rect -198 -62839 -94 -62441
rect 282 -62492 302 -62068
rect 366 -62492 386 -62068
rect 282 -62788 386 -62492
rect -307 -62840 15 -62839
rect -307 -63160 -306 -62840
rect 14 -63160 15 -62840
rect -307 -63161 15 -63160
rect -198 -63559 -94 -63161
rect 282 -63212 302 -62788
rect 366 -63212 386 -62788
rect 282 -63508 386 -63212
rect -307 -63560 15 -63559
rect -307 -63880 -306 -63560
rect 14 -63880 15 -63560
rect -307 -63881 15 -63880
rect -198 -64279 -94 -63881
rect 282 -63932 302 -63508
rect 366 -63932 386 -63508
rect 282 -64228 386 -63932
rect -307 -64280 15 -64279
rect -307 -64600 -306 -64280
rect 14 -64600 15 -64280
rect -307 -64601 15 -64600
rect -198 -64999 -94 -64601
rect 282 -64652 302 -64228
rect 366 -64652 386 -64228
rect 282 -64948 386 -64652
rect -307 -65000 15 -64999
rect -307 -65320 -306 -65000
rect 14 -65320 15 -65000
rect -307 -65321 15 -65320
rect -198 -65719 -94 -65321
rect 282 -65372 302 -64948
rect 366 -65372 386 -64948
rect 282 -65668 386 -65372
rect -307 -65720 15 -65719
rect -307 -66040 -306 -65720
rect 14 -66040 15 -65720
rect -307 -66041 15 -66040
rect -198 -66439 -94 -66041
rect 282 -66092 302 -65668
rect 366 -66092 386 -65668
rect 282 -66388 386 -66092
rect -307 -66440 15 -66439
rect -307 -66760 -306 -66440
rect 14 -66760 15 -66440
rect -307 -66761 15 -66760
rect -198 -67159 -94 -66761
rect 282 -66812 302 -66388
rect 366 -66812 386 -66388
rect 282 -67108 386 -66812
rect -307 -67160 15 -67159
rect -307 -67480 -306 -67160
rect 14 -67480 15 -67160
rect -307 -67481 15 -67480
rect -198 -67879 -94 -67481
rect 282 -67532 302 -67108
rect 366 -67532 386 -67108
rect 282 -67828 386 -67532
rect -307 -67880 15 -67879
rect -307 -68200 -306 -67880
rect 14 -68200 15 -67880
rect -307 -68201 15 -68200
rect -198 -68599 -94 -68201
rect 282 -68252 302 -67828
rect 366 -68252 386 -67828
rect 282 -68548 386 -68252
rect -307 -68600 15 -68599
rect -307 -68920 -306 -68600
rect 14 -68920 15 -68600
rect -307 -68921 15 -68920
rect -198 -69319 -94 -68921
rect 282 -68972 302 -68548
rect 366 -68972 386 -68548
rect 282 -69268 386 -68972
rect -307 -69320 15 -69319
rect -307 -69640 -306 -69320
rect 14 -69640 15 -69320
rect -307 -69641 15 -69640
rect -198 -70039 -94 -69641
rect 282 -69692 302 -69268
rect 366 -69692 386 -69268
rect 282 -69988 386 -69692
rect -307 -70040 15 -70039
rect -307 -70360 -306 -70040
rect 14 -70360 15 -70040
rect -307 -70361 15 -70360
rect -198 -70759 -94 -70361
rect 282 -70412 302 -69988
rect 366 -70412 386 -69988
rect 282 -70708 386 -70412
rect -307 -70760 15 -70759
rect -307 -71080 -306 -70760
rect 14 -71080 15 -70760
rect -307 -71081 15 -71080
rect -198 -71479 -94 -71081
rect 282 -71132 302 -70708
rect 366 -71132 386 -70708
rect 282 -71428 386 -71132
rect -307 -71480 15 -71479
rect -307 -71800 -306 -71480
rect 14 -71800 15 -71480
rect -307 -71801 15 -71800
rect -198 -72199 -94 -71801
rect 282 -71852 302 -71428
rect 366 -71852 386 -71428
rect 282 -72148 386 -71852
rect -307 -72200 15 -72199
rect -307 -72520 -306 -72200
rect 14 -72520 15 -72200
rect -307 -72521 15 -72520
rect -198 -72919 -94 -72521
rect 282 -72572 302 -72148
rect 366 -72572 386 -72148
rect 282 -72868 386 -72572
rect -307 -72920 15 -72919
rect -307 -73240 -306 -72920
rect 14 -73240 15 -72920
rect -307 -73241 15 -73240
rect -198 -73639 -94 -73241
rect 282 -73292 302 -72868
rect 366 -73292 386 -72868
rect 282 -73588 386 -73292
rect -307 -73640 15 -73639
rect -307 -73960 -306 -73640
rect 14 -73960 15 -73640
rect -307 -73961 15 -73960
rect -198 -74359 -94 -73961
rect 282 -74012 302 -73588
rect 366 -74012 386 -73588
rect 282 -74308 386 -74012
rect -307 -74360 15 -74359
rect -307 -74680 -306 -74360
rect 14 -74680 15 -74360
rect -307 -74681 15 -74680
rect -198 -75079 -94 -74681
rect 282 -74732 302 -74308
rect 366 -74732 386 -74308
rect 282 -75028 386 -74732
rect -307 -75080 15 -75079
rect -307 -75400 -306 -75080
rect 14 -75400 15 -75080
rect -307 -75401 15 -75400
rect -198 -75799 -94 -75401
rect 282 -75452 302 -75028
rect 366 -75452 386 -75028
rect 282 -75748 386 -75452
rect -307 -75800 15 -75799
rect -307 -76120 -306 -75800
rect 14 -76120 15 -75800
rect -307 -76121 15 -76120
rect -198 -76519 -94 -76121
rect 282 -76172 302 -75748
rect 366 -76172 386 -75748
rect 282 -76468 386 -76172
rect -307 -76520 15 -76519
rect -307 -76840 -306 -76520
rect 14 -76840 15 -76520
rect -307 -76841 15 -76840
rect -198 -77239 -94 -76841
rect 282 -76892 302 -76468
rect 366 -76892 386 -76468
rect 282 -77188 386 -76892
rect -307 -77240 15 -77239
rect -307 -77560 -306 -77240
rect 14 -77560 15 -77240
rect -307 -77561 15 -77560
rect -198 -77959 -94 -77561
rect 282 -77612 302 -77188
rect 366 -77612 386 -77188
rect 282 -77908 386 -77612
rect -307 -77960 15 -77959
rect -307 -78280 -306 -77960
rect 14 -78280 15 -77960
rect -307 -78281 15 -78280
rect -198 -78679 -94 -78281
rect 282 -78332 302 -77908
rect 366 -78332 386 -77908
rect 282 -78628 386 -78332
rect -307 -78680 15 -78679
rect -307 -79000 -306 -78680
rect 14 -79000 15 -78680
rect -307 -79001 15 -79000
rect -198 -79399 -94 -79001
rect 282 -79052 302 -78628
rect 366 -79052 386 -78628
rect 282 -79348 386 -79052
rect -307 -79400 15 -79399
rect -307 -79720 -306 -79400
rect 14 -79720 15 -79400
rect -307 -79721 15 -79720
rect -198 -80119 -94 -79721
rect 282 -79772 302 -79348
rect 366 -79772 386 -79348
rect 282 -80068 386 -79772
rect -307 -80120 15 -80119
rect -307 -80440 -306 -80120
rect 14 -80440 15 -80120
rect -307 -80441 15 -80440
rect -198 -80839 -94 -80441
rect 282 -80492 302 -80068
rect 366 -80492 386 -80068
rect 282 -80788 386 -80492
rect -307 -80840 15 -80839
rect -307 -81160 -306 -80840
rect 14 -81160 15 -80840
rect -307 -81161 15 -81160
rect -198 -81559 -94 -81161
rect 282 -81212 302 -80788
rect 366 -81212 386 -80788
rect 282 -81508 386 -81212
rect -307 -81560 15 -81559
rect -307 -81880 -306 -81560
rect 14 -81880 15 -81560
rect -307 -81881 15 -81880
rect -198 -82279 -94 -81881
rect 282 -81932 302 -81508
rect 366 -81932 386 -81508
rect 282 -82228 386 -81932
rect -307 -82280 15 -82279
rect -307 -82600 -306 -82280
rect 14 -82600 15 -82280
rect -307 -82601 15 -82600
rect -198 -82999 -94 -82601
rect 282 -82652 302 -82228
rect 366 -82652 386 -82228
rect 282 -82948 386 -82652
rect -307 -83000 15 -82999
rect -307 -83320 -306 -83000
rect 14 -83320 15 -83000
rect -307 -83321 15 -83320
rect -198 -83719 -94 -83321
rect 282 -83372 302 -82948
rect 366 -83372 386 -82948
rect 282 -83668 386 -83372
rect -307 -83720 15 -83719
rect -307 -84040 -306 -83720
rect 14 -84040 15 -83720
rect -307 -84041 15 -84040
rect -198 -84439 -94 -84041
rect 282 -84092 302 -83668
rect 366 -84092 386 -83668
rect 282 -84388 386 -84092
rect -307 -84440 15 -84439
rect -307 -84760 -306 -84440
rect 14 -84760 15 -84440
rect -307 -84761 15 -84760
rect -198 -85159 -94 -84761
rect 282 -84812 302 -84388
rect 366 -84812 386 -84388
rect 282 -85108 386 -84812
rect -307 -85160 15 -85159
rect -307 -85480 -306 -85160
rect 14 -85480 15 -85160
rect -307 -85481 15 -85480
rect -198 -85879 -94 -85481
rect 282 -85532 302 -85108
rect 366 -85532 386 -85108
rect 282 -85828 386 -85532
rect -307 -85880 15 -85879
rect -307 -86200 -306 -85880
rect 14 -86200 15 -85880
rect -307 -86201 15 -86200
rect -198 -86599 -94 -86201
rect 282 -86252 302 -85828
rect 366 -86252 386 -85828
rect 282 -86548 386 -86252
rect -307 -86600 15 -86599
rect -307 -86920 -306 -86600
rect 14 -86920 15 -86600
rect -307 -86921 15 -86920
rect -198 -87319 -94 -86921
rect 282 -86972 302 -86548
rect 366 -86972 386 -86548
rect 282 -87268 386 -86972
rect -307 -87320 15 -87319
rect -307 -87640 -306 -87320
rect 14 -87640 15 -87320
rect -307 -87641 15 -87640
rect -198 -88039 -94 -87641
rect 282 -87692 302 -87268
rect 366 -87692 386 -87268
rect 282 -87988 386 -87692
rect -307 -88040 15 -88039
rect -307 -88360 -306 -88040
rect 14 -88360 15 -88040
rect -307 -88361 15 -88360
rect -198 -88759 -94 -88361
rect 282 -88412 302 -87988
rect 366 -88412 386 -87988
rect 282 -88708 386 -88412
rect -307 -88760 15 -88759
rect -307 -89080 -306 -88760
rect 14 -89080 15 -88760
rect -307 -89081 15 -89080
rect -198 -89479 -94 -89081
rect 282 -89132 302 -88708
rect 366 -89132 386 -88708
rect 282 -89428 386 -89132
rect -307 -89480 15 -89479
rect -307 -89800 -306 -89480
rect 14 -89800 15 -89480
rect -307 -89801 15 -89800
rect -198 -90199 -94 -89801
rect 282 -89852 302 -89428
rect 366 -89852 386 -89428
rect 282 -90148 386 -89852
rect -307 -90200 15 -90199
rect -307 -90520 -306 -90200
rect 14 -90520 15 -90200
rect -307 -90521 15 -90520
rect -198 -90919 -94 -90521
rect 282 -90572 302 -90148
rect 366 -90572 386 -90148
rect 282 -90868 386 -90572
rect -307 -90920 15 -90919
rect -307 -91240 -306 -90920
rect 14 -91240 15 -90920
rect -307 -91241 15 -91240
rect -198 -91639 -94 -91241
rect 282 -91292 302 -90868
rect 366 -91292 386 -90868
rect 282 -91588 386 -91292
rect -307 -91640 15 -91639
rect -307 -91960 -306 -91640
rect 14 -91960 15 -91640
rect -307 -91961 15 -91960
rect -198 -92160 -94 -91961
rect 282 -92012 302 -91588
rect 366 -92012 386 -91588
rect 282 -92160 386 -92012
<< properties >>
string FIXED_BBOX -386 91560 94 92040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.0 l 2.0 val 9.52 carea 2.00 cperi 0.19 nx 1 ny 256 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
