magic
tech sky130A
timestamp 1728967704
<< nwell >>
rect -180 150 160 320
<< nmos >>
rect -5 -25 10 75
<< pmos >>
rect -5 180 10 280
<< ndiff >>
rect -55 55 -5 75
rect -55 -15 -45 55
rect -15 -15 -5 55
rect -55 -25 -5 -15
rect 10 55 75 75
rect 10 -15 30 55
rect 60 -15 75 55
rect 10 -25 75 -15
<< pdiff >>
rect -55 265 -5 280
rect -55 195 -45 265
rect -15 195 -5 265
rect -55 180 -5 195
rect 10 265 75 280
rect 10 195 30 265
rect 60 195 75 265
rect 10 180 75 195
<< ndiffc >>
rect -45 -15 -15 55
rect 30 -15 60 55
<< pdiffc >>
rect -45 195 -15 265
rect 30 195 60 265
<< psubdiff >>
rect -165 15 -100 30
rect -165 -30 -150 15
rect -115 -30 -100 15
rect -165 -45 -100 -30
<< nsubdiff >>
rect -150 255 -85 270
rect -150 210 -135 255
rect -100 210 -85 255
rect -150 185 -85 210
<< psubdiffcont >>
rect -150 -30 -115 15
<< nsubdiffcont >>
rect -135 210 -100 255
<< poly >>
rect -5 280 10 305
rect -5 125 10 180
rect -180 85 10 125
rect -5 75 10 85
rect -5 -40 10 -25
<< locali >>
rect -180 360 160 415
rect -150 255 -85 360
rect -150 210 -135 255
rect -100 210 -85 255
rect -150 185 -85 210
rect -50 265 -10 360
rect -50 195 -45 265
rect -15 195 -10 265
rect -50 185 -10 195
rect 20 265 70 280
rect 20 195 30 265
rect 60 195 70 265
rect 20 130 70 195
rect 20 85 160 130
rect -50 55 -10 65
rect -165 15 -100 30
rect -165 -30 -150 15
rect -115 -30 -100 15
rect -165 -90 -100 -30
rect -50 -15 -45 55
rect -15 -15 -10 55
rect -50 -90 -10 -15
rect 20 55 70 85
rect 20 -15 30 55
rect 60 -15 70 55
rect 20 -30 70 -15
rect -190 -145 165 -90
<< labels >>
rlabel locali 150 100 160 115 3 out
port 3 e
rlabel locali 150 -135 165 -120 3 gnd
port 4 e
rlabel locali 145 380 160 395 3 vdd
port 1 e
rlabel poly -180 95 -165 110 3 in
port 2 e
<< end >>
