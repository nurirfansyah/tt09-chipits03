magic
tech sky130A
magscale 1 2
timestamp 1730269323
<< metal3 >>
rect -386 5612 386 5640
rect -386 5188 302 5612
rect 366 5188 386 5612
rect -386 5160 386 5188
rect -386 4892 386 4920
rect -386 4468 302 4892
rect 366 4468 386 4892
rect -386 4440 386 4468
rect -386 4172 386 4200
rect -386 3748 302 4172
rect 366 3748 386 4172
rect -386 3720 386 3748
rect -386 3452 386 3480
rect -386 3028 302 3452
rect 366 3028 386 3452
rect -386 3000 386 3028
rect -386 2732 386 2760
rect -386 2308 302 2732
rect 366 2308 386 2732
rect -386 2280 386 2308
rect -386 2012 386 2040
rect -386 1588 302 2012
rect 366 1588 386 2012
rect -386 1560 386 1588
rect -386 1292 386 1320
rect -386 868 302 1292
rect 366 868 386 1292
rect -386 840 386 868
rect -386 572 386 600
rect -386 148 302 572
rect 366 148 386 572
rect -386 120 386 148
rect -386 -148 386 -120
rect -386 -572 302 -148
rect 366 -572 386 -148
rect -386 -600 386 -572
rect -386 -868 386 -840
rect -386 -1292 302 -868
rect 366 -1292 386 -868
rect -386 -1320 386 -1292
rect -386 -1588 386 -1560
rect -386 -2012 302 -1588
rect 366 -2012 386 -1588
rect -386 -2040 386 -2012
rect -386 -2308 386 -2280
rect -386 -2732 302 -2308
rect 366 -2732 386 -2308
rect -386 -2760 386 -2732
rect -386 -3028 386 -3000
rect -386 -3452 302 -3028
rect 366 -3452 386 -3028
rect -386 -3480 386 -3452
rect -386 -3748 386 -3720
rect -386 -4172 302 -3748
rect 366 -4172 386 -3748
rect -386 -4200 386 -4172
rect -386 -4468 386 -4440
rect -386 -4892 302 -4468
rect 366 -4892 386 -4468
rect -386 -4920 386 -4892
rect -386 -5188 386 -5160
rect -386 -5612 302 -5188
rect 366 -5612 386 -5188
rect -386 -5640 386 -5612
<< via3 >>
rect 302 5188 366 5612
rect 302 4468 366 4892
rect 302 3748 366 4172
rect 302 3028 366 3452
rect 302 2308 366 2732
rect 302 1588 366 2012
rect 302 868 366 1292
rect 302 148 366 572
rect 302 -572 366 -148
rect 302 -1292 366 -868
rect 302 -2012 366 -1588
rect 302 -2732 366 -2308
rect 302 -3452 366 -3028
rect 302 -4172 366 -3748
rect 302 -4892 366 -4468
rect 302 -5612 366 -5188
<< mimcap >>
rect -346 5560 54 5600
rect -346 5240 -306 5560
rect 14 5240 54 5560
rect -346 5200 54 5240
rect -346 4840 54 4880
rect -346 4520 -306 4840
rect 14 4520 54 4840
rect -346 4480 54 4520
rect -346 4120 54 4160
rect -346 3800 -306 4120
rect 14 3800 54 4120
rect -346 3760 54 3800
rect -346 3400 54 3440
rect -346 3080 -306 3400
rect 14 3080 54 3400
rect -346 3040 54 3080
rect -346 2680 54 2720
rect -346 2360 -306 2680
rect 14 2360 54 2680
rect -346 2320 54 2360
rect -346 1960 54 2000
rect -346 1640 -306 1960
rect 14 1640 54 1960
rect -346 1600 54 1640
rect -346 1240 54 1280
rect -346 920 -306 1240
rect 14 920 54 1240
rect -346 880 54 920
rect -346 520 54 560
rect -346 200 -306 520
rect 14 200 54 520
rect -346 160 54 200
rect -346 -200 54 -160
rect -346 -520 -306 -200
rect 14 -520 54 -200
rect -346 -560 54 -520
rect -346 -920 54 -880
rect -346 -1240 -306 -920
rect 14 -1240 54 -920
rect -346 -1280 54 -1240
rect -346 -1640 54 -1600
rect -346 -1960 -306 -1640
rect 14 -1960 54 -1640
rect -346 -2000 54 -1960
rect -346 -2360 54 -2320
rect -346 -2680 -306 -2360
rect 14 -2680 54 -2360
rect -346 -2720 54 -2680
rect -346 -3080 54 -3040
rect -346 -3400 -306 -3080
rect 14 -3400 54 -3080
rect -346 -3440 54 -3400
rect -346 -3800 54 -3760
rect -346 -4120 -306 -3800
rect 14 -4120 54 -3800
rect -346 -4160 54 -4120
rect -346 -4520 54 -4480
rect -346 -4840 -306 -4520
rect 14 -4840 54 -4520
rect -346 -4880 54 -4840
rect -346 -5240 54 -5200
rect -346 -5560 -306 -5240
rect 14 -5560 54 -5240
rect -346 -5600 54 -5560
<< mimcapcontact >>
rect -306 5240 14 5560
rect -306 4520 14 4840
rect -306 3800 14 4120
rect -306 3080 14 3400
rect -306 2360 14 2680
rect -306 1640 14 1960
rect -306 920 14 1240
rect -306 200 14 520
rect -306 -520 14 -200
rect -306 -1240 14 -920
rect -306 -1960 14 -1640
rect -306 -2680 14 -2360
rect -306 -3400 14 -3080
rect -306 -4120 14 -3800
rect -306 -4840 14 -4520
rect -306 -5560 14 -5240
<< metal4 >>
rect -198 5561 -94 5760
rect 282 5612 386 5760
rect -307 5560 15 5561
rect -307 5240 -306 5560
rect 14 5240 15 5560
rect -307 5239 15 5240
rect -198 4841 -94 5239
rect 282 5188 302 5612
rect 366 5188 386 5612
rect 282 4892 386 5188
rect -307 4840 15 4841
rect -307 4520 -306 4840
rect 14 4520 15 4840
rect -307 4519 15 4520
rect -198 4121 -94 4519
rect 282 4468 302 4892
rect 366 4468 386 4892
rect 282 4172 386 4468
rect -307 4120 15 4121
rect -307 3800 -306 4120
rect 14 3800 15 4120
rect -307 3799 15 3800
rect -198 3401 -94 3799
rect 282 3748 302 4172
rect 366 3748 386 4172
rect 282 3452 386 3748
rect -307 3400 15 3401
rect -307 3080 -306 3400
rect 14 3080 15 3400
rect -307 3079 15 3080
rect -198 2681 -94 3079
rect 282 3028 302 3452
rect 366 3028 386 3452
rect 282 2732 386 3028
rect -307 2680 15 2681
rect -307 2360 -306 2680
rect 14 2360 15 2680
rect -307 2359 15 2360
rect -198 1961 -94 2359
rect 282 2308 302 2732
rect 366 2308 386 2732
rect 282 2012 386 2308
rect -307 1960 15 1961
rect -307 1640 -306 1960
rect 14 1640 15 1960
rect -307 1639 15 1640
rect -198 1241 -94 1639
rect 282 1588 302 2012
rect 366 1588 386 2012
rect 282 1292 386 1588
rect -307 1240 15 1241
rect -307 920 -306 1240
rect 14 920 15 1240
rect -307 919 15 920
rect -198 521 -94 919
rect 282 868 302 1292
rect 366 868 386 1292
rect 282 572 386 868
rect -307 520 15 521
rect -307 200 -306 520
rect 14 200 15 520
rect -307 199 15 200
rect -198 -199 -94 199
rect 282 148 302 572
rect 366 148 386 572
rect 282 -148 386 148
rect -307 -200 15 -199
rect -307 -520 -306 -200
rect 14 -520 15 -200
rect -307 -521 15 -520
rect -198 -919 -94 -521
rect 282 -572 302 -148
rect 366 -572 386 -148
rect 282 -868 386 -572
rect -307 -920 15 -919
rect -307 -1240 -306 -920
rect 14 -1240 15 -920
rect -307 -1241 15 -1240
rect -198 -1639 -94 -1241
rect 282 -1292 302 -868
rect 366 -1292 386 -868
rect 282 -1588 386 -1292
rect -307 -1640 15 -1639
rect -307 -1960 -306 -1640
rect 14 -1960 15 -1640
rect -307 -1961 15 -1960
rect -198 -2359 -94 -1961
rect 282 -2012 302 -1588
rect 366 -2012 386 -1588
rect 282 -2308 386 -2012
rect -307 -2360 15 -2359
rect -307 -2680 -306 -2360
rect 14 -2680 15 -2360
rect -307 -2681 15 -2680
rect -198 -3079 -94 -2681
rect 282 -2732 302 -2308
rect 366 -2732 386 -2308
rect 282 -3028 386 -2732
rect -307 -3080 15 -3079
rect -307 -3400 -306 -3080
rect 14 -3400 15 -3080
rect -307 -3401 15 -3400
rect -198 -3799 -94 -3401
rect 282 -3452 302 -3028
rect 366 -3452 386 -3028
rect 282 -3748 386 -3452
rect -307 -3800 15 -3799
rect -307 -4120 -306 -3800
rect 14 -4120 15 -3800
rect -307 -4121 15 -4120
rect -198 -4519 -94 -4121
rect 282 -4172 302 -3748
rect 366 -4172 386 -3748
rect 282 -4468 386 -4172
rect -307 -4520 15 -4519
rect -307 -4840 -306 -4520
rect 14 -4840 15 -4520
rect -307 -4841 15 -4840
rect -198 -5239 -94 -4841
rect 282 -4892 302 -4468
rect 366 -4892 386 -4468
rect 282 -5188 386 -4892
rect -307 -5240 15 -5239
rect -307 -5560 -306 -5240
rect 14 -5560 15 -5240
rect -307 -5561 15 -5560
rect -198 -5760 -94 -5561
rect 282 -5612 302 -5188
rect 366 -5612 386 -5188
rect 282 -5760 386 -5612
<< properties >>
string FIXED_BBOX -386 5160 94 5640
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.0 l 2.0 val 9.52 carea 2.00 cperi 0.19 nx 1 ny 16 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
