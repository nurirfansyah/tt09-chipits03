magic
tech sky130A
magscale 1 2
timestamp 1730624594
<< metal3 >>
rect -7470 11372 -6698 11400
rect -7470 10948 -6782 11372
rect -6718 10948 -6698 11372
rect -7470 10920 -6698 10948
rect -6458 11372 -5686 11400
rect -6458 10948 -5770 11372
rect -5706 10948 -5686 11372
rect -6458 10920 -5686 10948
rect -5446 11372 -4674 11400
rect -5446 10948 -4758 11372
rect -4694 10948 -4674 11372
rect -5446 10920 -4674 10948
rect -4434 11372 -3662 11400
rect -4434 10948 -3746 11372
rect -3682 10948 -3662 11372
rect -4434 10920 -3662 10948
rect -3422 11372 -2650 11400
rect -3422 10948 -2734 11372
rect -2670 10948 -2650 11372
rect -3422 10920 -2650 10948
rect -2410 11372 -1638 11400
rect -2410 10948 -1722 11372
rect -1658 10948 -1638 11372
rect -2410 10920 -1638 10948
rect -1398 11372 -626 11400
rect -1398 10948 -710 11372
rect -646 10948 -626 11372
rect -1398 10920 -626 10948
rect -386 11372 386 11400
rect -386 10948 302 11372
rect 366 10948 386 11372
rect -386 10920 386 10948
rect 626 11372 1398 11400
rect 626 10948 1314 11372
rect 1378 10948 1398 11372
rect 626 10920 1398 10948
rect 1638 11372 2410 11400
rect 1638 10948 2326 11372
rect 2390 10948 2410 11372
rect 1638 10920 2410 10948
rect 2650 11372 3422 11400
rect 2650 10948 3338 11372
rect 3402 10948 3422 11372
rect 2650 10920 3422 10948
rect 3662 11372 4434 11400
rect 3662 10948 4350 11372
rect 4414 10948 4434 11372
rect 3662 10920 4434 10948
rect 4674 11372 5446 11400
rect 4674 10948 5362 11372
rect 5426 10948 5446 11372
rect 4674 10920 5446 10948
rect 5686 11372 6458 11400
rect 5686 10948 6374 11372
rect 6438 10948 6458 11372
rect 5686 10920 6458 10948
rect 6698 11372 7470 11400
rect 6698 10948 7386 11372
rect 7450 10948 7470 11372
rect 6698 10920 7470 10948
rect -7470 10652 -6698 10680
rect -7470 10228 -6782 10652
rect -6718 10228 -6698 10652
rect -7470 10200 -6698 10228
rect -6458 10652 -5686 10680
rect -6458 10228 -5770 10652
rect -5706 10228 -5686 10652
rect -6458 10200 -5686 10228
rect -5446 10652 -4674 10680
rect -5446 10228 -4758 10652
rect -4694 10228 -4674 10652
rect -5446 10200 -4674 10228
rect -4434 10652 -3662 10680
rect -4434 10228 -3746 10652
rect -3682 10228 -3662 10652
rect -4434 10200 -3662 10228
rect -3422 10652 -2650 10680
rect -3422 10228 -2734 10652
rect -2670 10228 -2650 10652
rect -3422 10200 -2650 10228
rect -2410 10652 -1638 10680
rect -2410 10228 -1722 10652
rect -1658 10228 -1638 10652
rect -2410 10200 -1638 10228
rect -1398 10652 -626 10680
rect -1398 10228 -710 10652
rect -646 10228 -626 10652
rect -1398 10200 -626 10228
rect -386 10652 386 10680
rect -386 10228 302 10652
rect 366 10228 386 10652
rect -386 10200 386 10228
rect 626 10652 1398 10680
rect 626 10228 1314 10652
rect 1378 10228 1398 10652
rect 626 10200 1398 10228
rect 1638 10652 2410 10680
rect 1638 10228 2326 10652
rect 2390 10228 2410 10652
rect 1638 10200 2410 10228
rect 2650 10652 3422 10680
rect 2650 10228 3338 10652
rect 3402 10228 3422 10652
rect 2650 10200 3422 10228
rect 3662 10652 4434 10680
rect 3662 10228 4350 10652
rect 4414 10228 4434 10652
rect 3662 10200 4434 10228
rect 4674 10652 5446 10680
rect 4674 10228 5362 10652
rect 5426 10228 5446 10652
rect 4674 10200 5446 10228
rect 5686 10652 6458 10680
rect 5686 10228 6374 10652
rect 6438 10228 6458 10652
rect 5686 10200 6458 10228
rect 6698 10652 7470 10680
rect 6698 10228 7386 10652
rect 7450 10228 7470 10652
rect 6698 10200 7470 10228
rect -7470 9932 -6698 9960
rect -7470 9508 -6782 9932
rect -6718 9508 -6698 9932
rect -7470 9480 -6698 9508
rect -6458 9932 -5686 9960
rect -6458 9508 -5770 9932
rect -5706 9508 -5686 9932
rect -6458 9480 -5686 9508
rect -5446 9932 -4674 9960
rect -5446 9508 -4758 9932
rect -4694 9508 -4674 9932
rect -5446 9480 -4674 9508
rect -4434 9932 -3662 9960
rect -4434 9508 -3746 9932
rect -3682 9508 -3662 9932
rect -4434 9480 -3662 9508
rect -3422 9932 -2650 9960
rect -3422 9508 -2734 9932
rect -2670 9508 -2650 9932
rect -3422 9480 -2650 9508
rect -2410 9932 -1638 9960
rect -2410 9508 -1722 9932
rect -1658 9508 -1638 9932
rect -2410 9480 -1638 9508
rect -1398 9932 -626 9960
rect -1398 9508 -710 9932
rect -646 9508 -626 9932
rect -1398 9480 -626 9508
rect -386 9932 386 9960
rect -386 9508 302 9932
rect 366 9508 386 9932
rect -386 9480 386 9508
rect 626 9932 1398 9960
rect 626 9508 1314 9932
rect 1378 9508 1398 9932
rect 626 9480 1398 9508
rect 1638 9932 2410 9960
rect 1638 9508 2326 9932
rect 2390 9508 2410 9932
rect 1638 9480 2410 9508
rect 2650 9932 3422 9960
rect 2650 9508 3338 9932
rect 3402 9508 3422 9932
rect 2650 9480 3422 9508
rect 3662 9932 4434 9960
rect 3662 9508 4350 9932
rect 4414 9508 4434 9932
rect 3662 9480 4434 9508
rect 4674 9932 5446 9960
rect 4674 9508 5362 9932
rect 5426 9508 5446 9932
rect 4674 9480 5446 9508
rect 5686 9932 6458 9960
rect 5686 9508 6374 9932
rect 6438 9508 6458 9932
rect 5686 9480 6458 9508
rect 6698 9932 7470 9960
rect 6698 9508 7386 9932
rect 7450 9508 7470 9932
rect 6698 9480 7470 9508
rect -7470 9212 -6698 9240
rect -7470 8788 -6782 9212
rect -6718 8788 -6698 9212
rect -7470 8760 -6698 8788
rect -6458 9212 -5686 9240
rect -6458 8788 -5770 9212
rect -5706 8788 -5686 9212
rect -6458 8760 -5686 8788
rect -5446 9212 -4674 9240
rect -5446 8788 -4758 9212
rect -4694 8788 -4674 9212
rect -5446 8760 -4674 8788
rect -4434 9212 -3662 9240
rect -4434 8788 -3746 9212
rect -3682 8788 -3662 9212
rect -4434 8760 -3662 8788
rect -3422 9212 -2650 9240
rect -3422 8788 -2734 9212
rect -2670 8788 -2650 9212
rect -3422 8760 -2650 8788
rect -2410 9212 -1638 9240
rect -2410 8788 -1722 9212
rect -1658 8788 -1638 9212
rect -2410 8760 -1638 8788
rect -1398 9212 -626 9240
rect -1398 8788 -710 9212
rect -646 8788 -626 9212
rect -1398 8760 -626 8788
rect -386 9212 386 9240
rect -386 8788 302 9212
rect 366 8788 386 9212
rect -386 8760 386 8788
rect 626 9212 1398 9240
rect 626 8788 1314 9212
rect 1378 8788 1398 9212
rect 626 8760 1398 8788
rect 1638 9212 2410 9240
rect 1638 8788 2326 9212
rect 2390 8788 2410 9212
rect 1638 8760 2410 8788
rect 2650 9212 3422 9240
rect 2650 8788 3338 9212
rect 3402 8788 3422 9212
rect 2650 8760 3422 8788
rect 3662 9212 4434 9240
rect 3662 8788 4350 9212
rect 4414 8788 4434 9212
rect 3662 8760 4434 8788
rect 4674 9212 5446 9240
rect 4674 8788 5362 9212
rect 5426 8788 5446 9212
rect 4674 8760 5446 8788
rect 5686 9212 6458 9240
rect 5686 8788 6374 9212
rect 6438 8788 6458 9212
rect 5686 8760 6458 8788
rect 6698 9212 7470 9240
rect 6698 8788 7386 9212
rect 7450 8788 7470 9212
rect 6698 8760 7470 8788
rect -7470 8492 -6698 8520
rect -7470 8068 -6782 8492
rect -6718 8068 -6698 8492
rect -7470 8040 -6698 8068
rect -6458 8492 -5686 8520
rect -6458 8068 -5770 8492
rect -5706 8068 -5686 8492
rect -6458 8040 -5686 8068
rect -5446 8492 -4674 8520
rect -5446 8068 -4758 8492
rect -4694 8068 -4674 8492
rect -5446 8040 -4674 8068
rect -4434 8492 -3662 8520
rect -4434 8068 -3746 8492
rect -3682 8068 -3662 8492
rect -4434 8040 -3662 8068
rect -3422 8492 -2650 8520
rect -3422 8068 -2734 8492
rect -2670 8068 -2650 8492
rect -3422 8040 -2650 8068
rect -2410 8492 -1638 8520
rect -2410 8068 -1722 8492
rect -1658 8068 -1638 8492
rect -2410 8040 -1638 8068
rect -1398 8492 -626 8520
rect -1398 8068 -710 8492
rect -646 8068 -626 8492
rect -1398 8040 -626 8068
rect -386 8492 386 8520
rect -386 8068 302 8492
rect 366 8068 386 8492
rect -386 8040 386 8068
rect 626 8492 1398 8520
rect 626 8068 1314 8492
rect 1378 8068 1398 8492
rect 626 8040 1398 8068
rect 1638 8492 2410 8520
rect 1638 8068 2326 8492
rect 2390 8068 2410 8492
rect 1638 8040 2410 8068
rect 2650 8492 3422 8520
rect 2650 8068 3338 8492
rect 3402 8068 3422 8492
rect 2650 8040 3422 8068
rect 3662 8492 4434 8520
rect 3662 8068 4350 8492
rect 4414 8068 4434 8492
rect 3662 8040 4434 8068
rect 4674 8492 5446 8520
rect 4674 8068 5362 8492
rect 5426 8068 5446 8492
rect 4674 8040 5446 8068
rect 5686 8492 6458 8520
rect 5686 8068 6374 8492
rect 6438 8068 6458 8492
rect 5686 8040 6458 8068
rect 6698 8492 7470 8520
rect 6698 8068 7386 8492
rect 7450 8068 7470 8492
rect 6698 8040 7470 8068
rect -7470 7772 -6698 7800
rect -7470 7348 -6782 7772
rect -6718 7348 -6698 7772
rect -7470 7320 -6698 7348
rect -6458 7772 -5686 7800
rect -6458 7348 -5770 7772
rect -5706 7348 -5686 7772
rect -6458 7320 -5686 7348
rect -5446 7772 -4674 7800
rect -5446 7348 -4758 7772
rect -4694 7348 -4674 7772
rect -5446 7320 -4674 7348
rect -4434 7772 -3662 7800
rect -4434 7348 -3746 7772
rect -3682 7348 -3662 7772
rect -4434 7320 -3662 7348
rect -3422 7772 -2650 7800
rect -3422 7348 -2734 7772
rect -2670 7348 -2650 7772
rect -3422 7320 -2650 7348
rect -2410 7772 -1638 7800
rect -2410 7348 -1722 7772
rect -1658 7348 -1638 7772
rect -2410 7320 -1638 7348
rect -1398 7772 -626 7800
rect -1398 7348 -710 7772
rect -646 7348 -626 7772
rect -1398 7320 -626 7348
rect -386 7772 386 7800
rect -386 7348 302 7772
rect 366 7348 386 7772
rect -386 7320 386 7348
rect 626 7772 1398 7800
rect 626 7348 1314 7772
rect 1378 7348 1398 7772
rect 626 7320 1398 7348
rect 1638 7772 2410 7800
rect 1638 7348 2326 7772
rect 2390 7348 2410 7772
rect 1638 7320 2410 7348
rect 2650 7772 3422 7800
rect 2650 7348 3338 7772
rect 3402 7348 3422 7772
rect 2650 7320 3422 7348
rect 3662 7772 4434 7800
rect 3662 7348 4350 7772
rect 4414 7348 4434 7772
rect 3662 7320 4434 7348
rect 4674 7772 5446 7800
rect 4674 7348 5362 7772
rect 5426 7348 5446 7772
rect 4674 7320 5446 7348
rect 5686 7772 6458 7800
rect 5686 7348 6374 7772
rect 6438 7348 6458 7772
rect 5686 7320 6458 7348
rect 6698 7772 7470 7800
rect 6698 7348 7386 7772
rect 7450 7348 7470 7772
rect 6698 7320 7470 7348
rect -7470 7052 -6698 7080
rect -7470 6628 -6782 7052
rect -6718 6628 -6698 7052
rect -7470 6600 -6698 6628
rect -6458 7052 -5686 7080
rect -6458 6628 -5770 7052
rect -5706 6628 -5686 7052
rect -6458 6600 -5686 6628
rect -5446 7052 -4674 7080
rect -5446 6628 -4758 7052
rect -4694 6628 -4674 7052
rect -5446 6600 -4674 6628
rect -4434 7052 -3662 7080
rect -4434 6628 -3746 7052
rect -3682 6628 -3662 7052
rect -4434 6600 -3662 6628
rect -3422 7052 -2650 7080
rect -3422 6628 -2734 7052
rect -2670 6628 -2650 7052
rect -3422 6600 -2650 6628
rect -2410 7052 -1638 7080
rect -2410 6628 -1722 7052
rect -1658 6628 -1638 7052
rect -2410 6600 -1638 6628
rect -1398 7052 -626 7080
rect -1398 6628 -710 7052
rect -646 6628 -626 7052
rect -1398 6600 -626 6628
rect -386 7052 386 7080
rect -386 6628 302 7052
rect 366 6628 386 7052
rect -386 6600 386 6628
rect 626 7052 1398 7080
rect 626 6628 1314 7052
rect 1378 6628 1398 7052
rect 626 6600 1398 6628
rect 1638 7052 2410 7080
rect 1638 6628 2326 7052
rect 2390 6628 2410 7052
rect 1638 6600 2410 6628
rect 2650 7052 3422 7080
rect 2650 6628 3338 7052
rect 3402 6628 3422 7052
rect 2650 6600 3422 6628
rect 3662 7052 4434 7080
rect 3662 6628 4350 7052
rect 4414 6628 4434 7052
rect 3662 6600 4434 6628
rect 4674 7052 5446 7080
rect 4674 6628 5362 7052
rect 5426 6628 5446 7052
rect 4674 6600 5446 6628
rect 5686 7052 6458 7080
rect 5686 6628 6374 7052
rect 6438 6628 6458 7052
rect 5686 6600 6458 6628
rect 6698 7052 7470 7080
rect 6698 6628 7386 7052
rect 7450 6628 7470 7052
rect 6698 6600 7470 6628
rect -7470 6332 -6698 6360
rect -7470 5908 -6782 6332
rect -6718 5908 -6698 6332
rect -7470 5880 -6698 5908
rect -6458 6332 -5686 6360
rect -6458 5908 -5770 6332
rect -5706 5908 -5686 6332
rect -6458 5880 -5686 5908
rect -5446 6332 -4674 6360
rect -5446 5908 -4758 6332
rect -4694 5908 -4674 6332
rect -5446 5880 -4674 5908
rect -4434 6332 -3662 6360
rect -4434 5908 -3746 6332
rect -3682 5908 -3662 6332
rect -4434 5880 -3662 5908
rect -3422 6332 -2650 6360
rect -3422 5908 -2734 6332
rect -2670 5908 -2650 6332
rect -3422 5880 -2650 5908
rect -2410 6332 -1638 6360
rect -2410 5908 -1722 6332
rect -1658 5908 -1638 6332
rect -2410 5880 -1638 5908
rect -1398 6332 -626 6360
rect -1398 5908 -710 6332
rect -646 5908 -626 6332
rect -1398 5880 -626 5908
rect -386 6332 386 6360
rect -386 5908 302 6332
rect 366 5908 386 6332
rect -386 5880 386 5908
rect 626 6332 1398 6360
rect 626 5908 1314 6332
rect 1378 5908 1398 6332
rect 626 5880 1398 5908
rect 1638 6332 2410 6360
rect 1638 5908 2326 6332
rect 2390 5908 2410 6332
rect 1638 5880 2410 5908
rect 2650 6332 3422 6360
rect 2650 5908 3338 6332
rect 3402 5908 3422 6332
rect 2650 5880 3422 5908
rect 3662 6332 4434 6360
rect 3662 5908 4350 6332
rect 4414 5908 4434 6332
rect 3662 5880 4434 5908
rect 4674 6332 5446 6360
rect 4674 5908 5362 6332
rect 5426 5908 5446 6332
rect 4674 5880 5446 5908
rect 5686 6332 6458 6360
rect 5686 5908 6374 6332
rect 6438 5908 6458 6332
rect 5686 5880 6458 5908
rect 6698 6332 7470 6360
rect 6698 5908 7386 6332
rect 7450 5908 7470 6332
rect 6698 5880 7470 5908
rect -7470 5612 -6698 5640
rect -7470 5188 -6782 5612
rect -6718 5188 -6698 5612
rect -7470 5160 -6698 5188
rect -6458 5612 -5686 5640
rect -6458 5188 -5770 5612
rect -5706 5188 -5686 5612
rect -6458 5160 -5686 5188
rect -5446 5612 -4674 5640
rect -5446 5188 -4758 5612
rect -4694 5188 -4674 5612
rect -5446 5160 -4674 5188
rect -4434 5612 -3662 5640
rect -4434 5188 -3746 5612
rect -3682 5188 -3662 5612
rect -4434 5160 -3662 5188
rect -3422 5612 -2650 5640
rect -3422 5188 -2734 5612
rect -2670 5188 -2650 5612
rect -3422 5160 -2650 5188
rect -2410 5612 -1638 5640
rect -2410 5188 -1722 5612
rect -1658 5188 -1638 5612
rect -2410 5160 -1638 5188
rect -1398 5612 -626 5640
rect -1398 5188 -710 5612
rect -646 5188 -626 5612
rect -1398 5160 -626 5188
rect -386 5612 386 5640
rect -386 5188 302 5612
rect 366 5188 386 5612
rect -386 5160 386 5188
rect 626 5612 1398 5640
rect 626 5188 1314 5612
rect 1378 5188 1398 5612
rect 626 5160 1398 5188
rect 1638 5612 2410 5640
rect 1638 5188 2326 5612
rect 2390 5188 2410 5612
rect 1638 5160 2410 5188
rect 2650 5612 3422 5640
rect 2650 5188 3338 5612
rect 3402 5188 3422 5612
rect 2650 5160 3422 5188
rect 3662 5612 4434 5640
rect 3662 5188 4350 5612
rect 4414 5188 4434 5612
rect 3662 5160 4434 5188
rect 4674 5612 5446 5640
rect 4674 5188 5362 5612
rect 5426 5188 5446 5612
rect 4674 5160 5446 5188
rect 5686 5612 6458 5640
rect 5686 5188 6374 5612
rect 6438 5188 6458 5612
rect 5686 5160 6458 5188
rect 6698 5612 7470 5640
rect 6698 5188 7386 5612
rect 7450 5188 7470 5612
rect 6698 5160 7470 5188
rect -7470 4892 -6698 4920
rect -7470 4468 -6782 4892
rect -6718 4468 -6698 4892
rect -7470 4440 -6698 4468
rect -6458 4892 -5686 4920
rect -6458 4468 -5770 4892
rect -5706 4468 -5686 4892
rect -6458 4440 -5686 4468
rect -5446 4892 -4674 4920
rect -5446 4468 -4758 4892
rect -4694 4468 -4674 4892
rect -5446 4440 -4674 4468
rect -4434 4892 -3662 4920
rect -4434 4468 -3746 4892
rect -3682 4468 -3662 4892
rect -4434 4440 -3662 4468
rect -3422 4892 -2650 4920
rect -3422 4468 -2734 4892
rect -2670 4468 -2650 4892
rect -3422 4440 -2650 4468
rect -2410 4892 -1638 4920
rect -2410 4468 -1722 4892
rect -1658 4468 -1638 4892
rect -2410 4440 -1638 4468
rect -1398 4892 -626 4920
rect -1398 4468 -710 4892
rect -646 4468 -626 4892
rect -1398 4440 -626 4468
rect -386 4892 386 4920
rect -386 4468 302 4892
rect 366 4468 386 4892
rect -386 4440 386 4468
rect 626 4892 1398 4920
rect 626 4468 1314 4892
rect 1378 4468 1398 4892
rect 626 4440 1398 4468
rect 1638 4892 2410 4920
rect 1638 4468 2326 4892
rect 2390 4468 2410 4892
rect 1638 4440 2410 4468
rect 2650 4892 3422 4920
rect 2650 4468 3338 4892
rect 3402 4468 3422 4892
rect 2650 4440 3422 4468
rect 3662 4892 4434 4920
rect 3662 4468 4350 4892
rect 4414 4468 4434 4892
rect 3662 4440 4434 4468
rect 4674 4892 5446 4920
rect 4674 4468 5362 4892
rect 5426 4468 5446 4892
rect 4674 4440 5446 4468
rect 5686 4892 6458 4920
rect 5686 4468 6374 4892
rect 6438 4468 6458 4892
rect 5686 4440 6458 4468
rect 6698 4892 7470 4920
rect 6698 4468 7386 4892
rect 7450 4468 7470 4892
rect 6698 4440 7470 4468
rect -7470 4172 -6698 4200
rect -7470 3748 -6782 4172
rect -6718 3748 -6698 4172
rect -7470 3720 -6698 3748
rect -6458 4172 -5686 4200
rect -6458 3748 -5770 4172
rect -5706 3748 -5686 4172
rect -6458 3720 -5686 3748
rect -5446 4172 -4674 4200
rect -5446 3748 -4758 4172
rect -4694 3748 -4674 4172
rect -5446 3720 -4674 3748
rect -4434 4172 -3662 4200
rect -4434 3748 -3746 4172
rect -3682 3748 -3662 4172
rect -4434 3720 -3662 3748
rect -3422 4172 -2650 4200
rect -3422 3748 -2734 4172
rect -2670 3748 -2650 4172
rect -3422 3720 -2650 3748
rect -2410 4172 -1638 4200
rect -2410 3748 -1722 4172
rect -1658 3748 -1638 4172
rect -2410 3720 -1638 3748
rect -1398 4172 -626 4200
rect -1398 3748 -710 4172
rect -646 3748 -626 4172
rect -1398 3720 -626 3748
rect -386 4172 386 4200
rect -386 3748 302 4172
rect 366 3748 386 4172
rect -386 3720 386 3748
rect 626 4172 1398 4200
rect 626 3748 1314 4172
rect 1378 3748 1398 4172
rect 626 3720 1398 3748
rect 1638 4172 2410 4200
rect 1638 3748 2326 4172
rect 2390 3748 2410 4172
rect 1638 3720 2410 3748
rect 2650 4172 3422 4200
rect 2650 3748 3338 4172
rect 3402 3748 3422 4172
rect 2650 3720 3422 3748
rect 3662 4172 4434 4200
rect 3662 3748 4350 4172
rect 4414 3748 4434 4172
rect 3662 3720 4434 3748
rect 4674 4172 5446 4200
rect 4674 3748 5362 4172
rect 5426 3748 5446 4172
rect 4674 3720 5446 3748
rect 5686 4172 6458 4200
rect 5686 3748 6374 4172
rect 6438 3748 6458 4172
rect 5686 3720 6458 3748
rect 6698 4172 7470 4200
rect 6698 3748 7386 4172
rect 7450 3748 7470 4172
rect 6698 3720 7470 3748
rect -7470 3452 -6698 3480
rect -7470 3028 -6782 3452
rect -6718 3028 -6698 3452
rect -7470 3000 -6698 3028
rect -6458 3452 -5686 3480
rect -6458 3028 -5770 3452
rect -5706 3028 -5686 3452
rect -6458 3000 -5686 3028
rect -5446 3452 -4674 3480
rect -5446 3028 -4758 3452
rect -4694 3028 -4674 3452
rect -5446 3000 -4674 3028
rect -4434 3452 -3662 3480
rect -4434 3028 -3746 3452
rect -3682 3028 -3662 3452
rect -4434 3000 -3662 3028
rect -3422 3452 -2650 3480
rect -3422 3028 -2734 3452
rect -2670 3028 -2650 3452
rect -3422 3000 -2650 3028
rect -2410 3452 -1638 3480
rect -2410 3028 -1722 3452
rect -1658 3028 -1638 3452
rect -2410 3000 -1638 3028
rect -1398 3452 -626 3480
rect -1398 3028 -710 3452
rect -646 3028 -626 3452
rect -1398 3000 -626 3028
rect -386 3452 386 3480
rect -386 3028 302 3452
rect 366 3028 386 3452
rect -386 3000 386 3028
rect 626 3452 1398 3480
rect 626 3028 1314 3452
rect 1378 3028 1398 3452
rect 626 3000 1398 3028
rect 1638 3452 2410 3480
rect 1638 3028 2326 3452
rect 2390 3028 2410 3452
rect 1638 3000 2410 3028
rect 2650 3452 3422 3480
rect 2650 3028 3338 3452
rect 3402 3028 3422 3452
rect 2650 3000 3422 3028
rect 3662 3452 4434 3480
rect 3662 3028 4350 3452
rect 4414 3028 4434 3452
rect 3662 3000 4434 3028
rect 4674 3452 5446 3480
rect 4674 3028 5362 3452
rect 5426 3028 5446 3452
rect 4674 3000 5446 3028
rect 5686 3452 6458 3480
rect 5686 3028 6374 3452
rect 6438 3028 6458 3452
rect 5686 3000 6458 3028
rect 6698 3452 7470 3480
rect 6698 3028 7386 3452
rect 7450 3028 7470 3452
rect 6698 3000 7470 3028
rect -7470 2732 -6698 2760
rect -7470 2308 -6782 2732
rect -6718 2308 -6698 2732
rect -7470 2280 -6698 2308
rect -6458 2732 -5686 2760
rect -6458 2308 -5770 2732
rect -5706 2308 -5686 2732
rect -6458 2280 -5686 2308
rect -5446 2732 -4674 2760
rect -5446 2308 -4758 2732
rect -4694 2308 -4674 2732
rect -5446 2280 -4674 2308
rect -4434 2732 -3662 2760
rect -4434 2308 -3746 2732
rect -3682 2308 -3662 2732
rect -4434 2280 -3662 2308
rect -3422 2732 -2650 2760
rect -3422 2308 -2734 2732
rect -2670 2308 -2650 2732
rect -3422 2280 -2650 2308
rect -2410 2732 -1638 2760
rect -2410 2308 -1722 2732
rect -1658 2308 -1638 2732
rect -2410 2280 -1638 2308
rect -1398 2732 -626 2760
rect -1398 2308 -710 2732
rect -646 2308 -626 2732
rect -1398 2280 -626 2308
rect -386 2732 386 2760
rect -386 2308 302 2732
rect 366 2308 386 2732
rect -386 2280 386 2308
rect 626 2732 1398 2760
rect 626 2308 1314 2732
rect 1378 2308 1398 2732
rect 626 2280 1398 2308
rect 1638 2732 2410 2760
rect 1638 2308 2326 2732
rect 2390 2308 2410 2732
rect 1638 2280 2410 2308
rect 2650 2732 3422 2760
rect 2650 2308 3338 2732
rect 3402 2308 3422 2732
rect 2650 2280 3422 2308
rect 3662 2732 4434 2760
rect 3662 2308 4350 2732
rect 4414 2308 4434 2732
rect 3662 2280 4434 2308
rect 4674 2732 5446 2760
rect 4674 2308 5362 2732
rect 5426 2308 5446 2732
rect 4674 2280 5446 2308
rect 5686 2732 6458 2760
rect 5686 2308 6374 2732
rect 6438 2308 6458 2732
rect 5686 2280 6458 2308
rect 6698 2732 7470 2760
rect 6698 2308 7386 2732
rect 7450 2308 7470 2732
rect 6698 2280 7470 2308
rect -7470 2012 -6698 2040
rect -7470 1588 -6782 2012
rect -6718 1588 -6698 2012
rect -7470 1560 -6698 1588
rect -6458 2012 -5686 2040
rect -6458 1588 -5770 2012
rect -5706 1588 -5686 2012
rect -6458 1560 -5686 1588
rect -5446 2012 -4674 2040
rect -5446 1588 -4758 2012
rect -4694 1588 -4674 2012
rect -5446 1560 -4674 1588
rect -4434 2012 -3662 2040
rect -4434 1588 -3746 2012
rect -3682 1588 -3662 2012
rect -4434 1560 -3662 1588
rect -3422 2012 -2650 2040
rect -3422 1588 -2734 2012
rect -2670 1588 -2650 2012
rect -3422 1560 -2650 1588
rect -2410 2012 -1638 2040
rect -2410 1588 -1722 2012
rect -1658 1588 -1638 2012
rect -2410 1560 -1638 1588
rect -1398 2012 -626 2040
rect -1398 1588 -710 2012
rect -646 1588 -626 2012
rect -1398 1560 -626 1588
rect -386 2012 386 2040
rect -386 1588 302 2012
rect 366 1588 386 2012
rect -386 1560 386 1588
rect 626 2012 1398 2040
rect 626 1588 1314 2012
rect 1378 1588 1398 2012
rect 626 1560 1398 1588
rect 1638 2012 2410 2040
rect 1638 1588 2326 2012
rect 2390 1588 2410 2012
rect 1638 1560 2410 1588
rect 2650 2012 3422 2040
rect 2650 1588 3338 2012
rect 3402 1588 3422 2012
rect 2650 1560 3422 1588
rect 3662 2012 4434 2040
rect 3662 1588 4350 2012
rect 4414 1588 4434 2012
rect 3662 1560 4434 1588
rect 4674 2012 5446 2040
rect 4674 1588 5362 2012
rect 5426 1588 5446 2012
rect 4674 1560 5446 1588
rect 5686 2012 6458 2040
rect 5686 1588 6374 2012
rect 6438 1588 6458 2012
rect 5686 1560 6458 1588
rect 6698 2012 7470 2040
rect 6698 1588 7386 2012
rect 7450 1588 7470 2012
rect 6698 1560 7470 1588
rect -7470 1292 -6698 1320
rect -7470 868 -6782 1292
rect -6718 868 -6698 1292
rect -7470 840 -6698 868
rect -6458 1292 -5686 1320
rect -6458 868 -5770 1292
rect -5706 868 -5686 1292
rect -6458 840 -5686 868
rect -5446 1292 -4674 1320
rect -5446 868 -4758 1292
rect -4694 868 -4674 1292
rect -5446 840 -4674 868
rect -4434 1292 -3662 1320
rect -4434 868 -3746 1292
rect -3682 868 -3662 1292
rect -4434 840 -3662 868
rect -3422 1292 -2650 1320
rect -3422 868 -2734 1292
rect -2670 868 -2650 1292
rect -3422 840 -2650 868
rect -2410 1292 -1638 1320
rect -2410 868 -1722 1292
rect -1658 868 -1638 1292
rect -2410 840 -1638 868
rect -1398 1292 -626 1320
rect -1398 868 -710 1292
rect -646 868 -626 1292
rect -1398 840 -626 868
rect -386 1292 386 1320
rect -386 868 302 1292
rect 366 868 386 1292
rect -386 840 386 868
rect 626 1292 1398 1320
rect 626 868 1314 1292
rect 1378 868 1398 1292
rect 626 840 1398 868
rect 1638 1292 2410 1320
rect 1638 868 2326 1292
rect 2390 868 2410 1292
rect 1638 840 2410 868
rect 2650 1292 3422 1320
rect 2650 868 3338 1292
rect 3402 868 3422 1292
rect 2650 840 3422 868
rect 3662 1292 4434 1320
rect 3662 868 4350 1292
rect 4414 868 4434 1292
rect 3662 840 4434 868
rect 4674 1292 5446 1320
rect 4674 868 5362 1292
rect 5426 868 5446 1292
rect 4674 840 5446 868
rect 5686 1292 6458 1320
rect 5686 868 6374 1292
rect 6438 868 6458 1292
rect 5686 840 6458 868
rect 6698 1292 7470 1320
rect 6698 868 7386 1292
rect 7450 868 7470 1292
rect 6698 840 7470 868
rect -7470 572 -6698 600
rect -7470 148 -6782 572
rect -6718 148 -6698 572
rect -7470 120 -6698 148
rect -6458 572 -5686 600
rect -6458 148 -5770 572
rect -5706 148 -5686 572
rect -6458 120 -5686 148
rect -5446 572 -4674 600
rect -5446 148 -4758 572
rect -4694 148 -4674 572
rect -5446 120 -4674 148
rect -4434 572 -3662 600
rect -4434 148 -3746 572
rect -3682 148 -3662 572
rect -4434 120 -3662 148
rect -3422 572 -2650 600
rect -3422 148 -2734 572
rect -2670 148 -2650 572
rect -3422 120 -2650 148
rect -2410 572 -1638 600
rect -2410 148 -1722 572
rect -1658 148 -1638 572
rect -2410 120 -1638 148
rect -1398 572 -626 600
rect -1398 148 -710 572
rect -646 148 -626 572
rect -1398 120 -626 148
rect -386 572 386 600
rect -386 148 302 572
rect 366 148 386 572
rect -386 120 386 148
rect 626 572 1398 600
rect 626 148 1314 572
rect 1378 148 1398 572
rect 626 120 1398 148
rect 1638 572 2410 600
rect 1638 148 2326 572
rect 2390 148 2410 572
rect 1638 120 2410 148
rect 2650 572 3422 600
rect 2650 148 3338 572
rect 3402 148 3422 572
rect 2650 120 3422 148
rect 3662 572 4434 600
rect 3662 148 4350 572
rect 4414 148 4434 572
rect 3662 120 4434 148
rect 4674 572 5446 600
rect 4674 148 5362 572
rect 5426 148 5446 572
rect 4674 120 5446 148
rect 5686 572 6458 600
rect 5686 148 6374 572
rect 6438 148 6458 572
rect 5686 120 6458 148
rect 6698 572 7470 600
rect 6698 148 7386 572
rect 7450 148 7470 572
rect 6698 120 7470 148
rect -7470 -148 -6698 -120
rect -7470 -572 -6782 -148
rect -6718 -572 -6698 -148
rect -7470 -600 -6698 -572
rect -6458 -148 -5686 -120
rect -6458 -572 -5770 -148
rect -5706 -572 -5686 -148
rect -6458 -600 -5686 -572
rect -5446 -148 -4674 -120
rect -5446 -572 -4758 -148
rect -4694 -572 -4674 -148
rect -5446 -600 -4674 -572
rect -4434 -148 -3662 -120
rect -4434 -572 -3746 -148
rect -3682 -572 -3662 -148
rect -4434 -600 -3662 -572
rect -3422 -148 -2650 -120
rect -3422 -572 -2734 -148
rect -2670 -572 -2650 -148
rect -3422 -600 -2650 -572
rect -2410 -148 -1638 -120
rect -2410 -572 -1722 -148
rect -1658 -572 -1638 -148
rect -2410 -600 -1638 -572
rect -1398 -148 -626 -120
rect -1398 -572 -710 -148
rect -646 -572 -626 -148
rect -1398 -600 -626 -572
rect -386 -148 386 -120
rect -386 -572 302 -148
rect 366 -572 386 -148
rect -386 -600 386 -572
rect 626 -148 1398 -120
rect 626 -572 1314 -148
rect 1378 -572 1398 -148
rect 626 -600 1398 -572
rect 1638 -148 2410 -120
rect 1638 -572 2326 -148
rect 2390 -572 2410 -148
rect 1638 -600 2410 -572
rect 2650 -148 3422 -120
rect 2650 -572 3338 -148
rect 3402 -572 3422 -148
rect 2650 -600 3422 -572
rect 3662 -148 4434 -120
rect 3662 -572 4350 -148
rect 4414 -572 4434 -148
rect 3662 -600 4434 -572
rect 4674 -148 5446 -120
rect 4674 -572 5362 -148
rect 5426 -572 5446 -148
rect 4674 -600 5446 -572
rect 5686 -148 6458 -120
rect 5686 -572 6374 -148
rect 6438 -572 6458 -148
rect 5686 -600 6458 -572
rect 6698 -148 7470 -120
rect 6698 -572 7386 -148
rect 7450 -572 7470 -148
rect 6698 -600 7470 -572
rect -7470 -868 -6698 -840
rect -7470 -1292 -6782 -868
rect -6718 -1292 -6698 -868
rect -7470 -1320 -6698 -1292
rect -6458 -868 -5686 -840
rect -6458 -1292 -5770 -868
rect -5706 -1292 -5686 -868
rect -6458 -1320 -5686 -1292
rect -5446 -868 -4674 -840
rect -5446 -1292 -4758 -868
rect -4694 -1292 -4674 -868
rect -5446 -1320 -4674 -1292
rect -4434 -868 -3662 -840
rect -4434 -1292 -3746 -868
rect -3682 -1292 -3662 -868
rect -4434 -1320 -3662 -1292
rect -3422 -868 -2650 -840
rect -3422 -1292 -2734 -868
rect -2670 -1292 -2650 -868
rect -3422 -1320 -2650 -1292
rect -2410 -868 -1638 -840
rect -2410 -1292 -1722 -868
rect -1658 -1292 -1638 -868
rect -2410 -1320 -1638 -1292
rect -1398 -868 -626 -840
rect -1398 -1292 -710 -868
rect -646 -1292 -626 -868
rect -1398 -1320 -626 -1292
rect -386 -868 386 -840
rect -386 -1292 302 -868
rect 366 -1292 386 -868
rect -386 -1320 386 -1292
rect 626 -868 1398 -840
rect 626 -1292 1314 -868
rect 1378 -1292 1398 -868
rect 626 -1320 1398 -1292
rect 1638 -868 2410 -840
rect 1638 -1292 2326 -868
rect 2390 -1292 2410 -868
rect 1638 -1320 2410 -1292
rect 2650 -868 3422 -840
rect 2650 -1292 3338 -868
rect 3402 -1292 3422 -868
rect 2650 -1320 3422 -1292
rect 3662 -868 4434 -840
rect 3662 -1292 4350 -868
rect 4414 -1292 4434 -868
rect 3662 -1320 4434 -1292
rect 4674 -868 5446 -840
rect 4674 -1292 5362 -868
rect 5426 -1292 5446 -868
rect 4674 -1320 5446 -1292
rect 5686 -868 6458 -840
rect 5686 -1292 6374 -868
rect 6438 -1292 6458 -868
rect 5686 -1320 6458 -1292
rect 6698 -868 7470 -840
rect 6698 -1292 7386 -868
rect 7450 -1292 7470 -868
rect 6698 -1320 7470 -1292
rect -7470 -1588 -6698 -1560
rect -7470 -2012 -6782 -1588
rect -6718 -2012 -6698 -1588
rect -7470 -2040 -6698 -2012
rect -6458 -1588 -5686 -1560
rect -6458 -2012 -5770 -1588
rect -5706 -2012 -5686 -1588
rect -6458 -2040 -5686 -2012
rect -5446 -1588 -4674 -1560
rect -5446 -2012 -4758 -1588
rect -4694 -2012 -4674 -1588
rect -5446 -2040 -4674 -2012
rect -4434 -1588 -3662 -1560
rect -4434 -2012 -3746 -1588
rect -3682 -2012 -3662 -1588
rect -4434 -2040 -3662 -2012
rect -3422 -1588 -2650 -1560
rect -3422 -2012 -2734 -1588
rect -2670 -2012 -2650 -1588
rect -3422 -2040 -2650 -2012
rect -2410 -1588 -1638 -1560
rect -2410 -2012 -1722 -1588
rect -1658 -2012 -1638 -1588
rect -2410 -2040 -1638 -2012
rect -1398 -1588 -626 -1560
rect -1398 -2012 -710 -1588
rect -646 -2012 -626 -1588
rect -1398 -2040 -626 -2012
rect -386 -1588 386 -1560
rect -386 -2012 302 -1588
rect 366 -2012 386 -1588
rect -386 -2040 386 -2012
rect 626 -1588 1398 -1560
rect 626 -2012 1314 -1588
rect 1378 -2012 1398 -1588
rect 626 -2040 1398 -2012
rect 1638 -1588 2410 -1560
rect 1638 -2012 2326 -1588
rect 2390 -2012 2410 -1588
rect 1638 -2040 2410 -2012
rect 2650 -1588 3422 -1560
rect 2650 -2012 3338 -1588
rect 3402 -2012 3422 -1588
rect 2650 -2040 3422 -2012
rect 3662 -1588 4434 -1560
rect 3662 -2012 4350 -1588
rect 4414 -2012 4434 -1588
rect 3662 -2040 4434 -2012
rect 4674 -1588 5446 -1560
rect 4674 -2012 5362 -1588
rect 5426 -2012 5446 -1588
rect 4674 -2040 5446 -2012
rect 5686 -1588 6458 -1560
rect 5686 -2012 6374 -1588
rect 6438 -2012 6458 -1588
rect 5686 -2040 6458 -2012
rect 6698 -1588 7470 -1560
rect 6698 -2012 7386 -1588
rect 7450 -2012 7470 -1588
rect 6698 -2040 7470 -2012
rect -7470 -2308 -6698 -2280
rect -7470 -2732 -6782 -2308
rect -6718 -2732 -6698 -2308
rect -7470 -2760 -6698 -2732
rect -6458 -2308 -5686 -2280
rect -6458 -2732 -5770 -2308
rect -5706 -2732 -5686 -2308
rect -6458 -2760 -5686 -2732
rect -5446 -2308 -4674 -2280
rect -5446 -2732 -4758 -2308
rect -4694 -2732 -4674 -2308
rect -5446 -2760 -4674 -2732
rect -4434 -2308 -3662 -2280
rect -4434 -2732 -3746 -2308
rect -3682 -2732 -3662 -2308
rect -4434 -2760 -3662 -2732
rect -3422 -2308 -2650 -2280
rect -3422 -2732 -2734 -2308
rect -2670 -2732 -2650 -2308
rect -3422 -2760 -2650 -2732
rect -2410 -2308 -1638 -2280
rect -2410 -2732 -1722 -2308
rect -1658 -2732 -1638 -2308
rect -2410 -2760 -1638 -2732
rect -1398 -2308 -626 -2280
rect -1398 -2732 -710 -2308
rect -646 -2732 -626 -2308
rect -1398 -2760 -626 -2732
rect -386 -2308 386 -2280
rect -386 -2732 302 -2308
rect 366 -2732 386 -2308
rect -386 -2760 386 -2732
rect 626 -2308 1398 -2280
rect 626 -2732 1314 -2308
rect 1378 -2732 1398 -2308
rect 626 -2760 1398 -2732
rect 1638 -2308 2410 -2280
rect 1638 -2732 2326 -2308
rect 2390 -2732 2410 -2308
rect 1638 -2760 2410 -2732
rect 2650 -2308 3422 -2280
rect 2650 -2732 3338 -2308
rect 3402 -2732 3422 -2308
rect 2650 -2760 3422 -2732
rect 3662 -2308 4434 -2280
rect 3662 -2732 4350 -2308
rect 4414 -2732 4434 -2308
rect 3662 -2760 4434 -2732
rect 4674 -2308 5446 -2280
rect 4674 -2732 5362 -2308
rect 5426 -2732 5446 -2308
rect 4674 -2760 5446 -2732
rect 5686 -2308 6458 -2280
rect 5686 -2732 6374 -2308
rect 6438 -2732 6458 -2308
rect 5686 -2760 6458 -2732
rect 6698 -2308 7470 -2280
rect 6698 -2732 7386 -2308
rect 7450 -2732 7470 -2308
rect 6698 -2760 7470 -2732
rect -7470 -3028 -6698 -3000
rect -7470 -3452 -6782 -3028
rect -6718 -3452 -6698 -3028
rect -7470 -3480 -6698 -3452
rect -6458 -3028 -5686 -3000
rect -6458 -3452 -5770 -3028
rect -5706 -3452 -5686 -3028
rect -6458 -3480 -5686 -3452
rect -5446 -3028 -4674 -3000
rect -5446 -3452 -4758 -3028
rect -4694 -3452 -4674 -3028
rect -5446 -3480 -4674 -3452
rect -4434 -3028 -3662 -3000
rect -4434 -3452 -3746 -3028
rect -3682 -3452 -3662 -3028
rect -4434 -3480 -3662 -3452
rect -3422 -3028 -2650 -3000
rect -3422 -3452 -2734 -3028
rect -2670 -3452 -2650 -3028
rect -3422 -3480 -2650 -3452
rect -2410 -3028 -1638 -3000
rect -2410 -3452 -1722 -3028
rect -1658 -3452 -1638 -3028
rect -2410 -3480 -1638 -3452
rect -1398 -3028 -626 -3000
rect -1398 -3452 -710 -3028
rect -646 -3452 -626 -3028
rect -1398 -3480 -626 -3452
rect -386 -3028 386 -3000
rect -386 -3452 302 -3028
rect 366 -3452 386 -3028
rect -386 -3480 386 -3452
rect 626 -3028 1398 -3000
rect 626 -3452 1314 -3028
rect 1378 -3452 1398 -3028
rect 626 -3480 1398 -3452
rect 1638 -3028 2410 -3000
rect 1638 -3452 2326 -3028
rect 2390 -3452 2410 -3028
rect 1638 -3480 2410 -3452
rect 2650 -3028 3422 -3000
rect 2650 -3452 3338 -3028
rect 3402 -3452 3422 -3028
rect 2650 -3480 3422 -3452
rect 3662 -3028 4434 -3000
rect 3662 -3452 4350 -3028
rect 4414 -3452 4434 -3028
rect 3662 -3480 4434 -3452
rect 4674 -3028 5446 -3000
rect 4674 -3452 5362 -3028
rect 5426 -3452 5446 -3028
rect 4674 -3480 5446 -3452
rect 5686 -3028 6458 -3000
rect 5686 -3452 6374 -3028
rect 6438 -3452 6458 -3028
rect 5686 -3480 6458 -3452
rect 6698 -3028 7470 -3000
rect 6698 -3452 7386 -3028
rect 7450 -3452 7470 -3028
rect 6698 -3480 7470 -3452
rect -7470 -3748 -6698 -3720
rect -7470 -4172 -6782 -3748
rect -6718 -4172 -6698 -3748
rect -7470 -4200 -6698 -4172
rect -6458 -3748 -5686 -3720
rect -6458 -4172 -5770 -3748
rect -5706 -4172 -5686 -3748
rect -6458 -4200 -5686 -4172
rect -5446 -3748 -4674 -3720
rect -5446 -4172 -4758 -3748
rect -4694 -4172 -4674 -3748
rect -5446 -4200 -4674 -4172
rect -4434 -3748 -3662 -3720
rect -4434 -4172 -3746 -3748
rect -3682 -4172 -3662 -3748
rect -4434 -4200 -3662 -4172
rect -3422 -3748 -2650 -3720
rect -3422 -4172 -2734 -3748
rect -2670 -4172 -2650 -3748
rect -3422 -4200 -2650 -4172
rect -2410 -3748 -1638 -3720
rect -2410 -4172 -1722 -3748
rect -1658 -4172 -1638 -3748
rect -2410 -4200 -1638 -4172
rect -1398 -3748 -626 -3720
rect -1398 -4172 -710 -3748
rect -646 -4172 -626 -3748
rect -1398 -4200 -626 -4172
rect -386 -3748 386 -3720
rect -386 -4172 302 -3748
rect 366 -4172 386 -3748
rect -386 -4200 386 -4172
rect 626 -3748 1398 -3720
rect 626 -4172 1314 -3748
rect 1378 -4172 1398 -3748
rect 626 -4200 1398 -4172
rect 1638 -3748 2410 -3720
rect 1638 -4172 2326 -3748
rect 2390 -4172 2410 -3748
rect 1638 -4200 2410 -4172
rect 2650 -3748 3422 -3720
rect 2650 -4172 3338 -3748
rect 3402 -4172 3422 -3748
rect 2650 -4200 3422 -4172
rect 3662 -3748 4434 -3720
rect 3662 -4172 4350 -3748
rect 4414 -4172 4434 -3748
rect 3662 -4200 4434 -4172
rect 4674 -3748 5446 -3720
rect 4674 -4172 5362 -3748
rect 5426 -4172 5446 -3748
rect 4674 -4200 5446 -4172
rect 5686 -3748 6458 -3720
rect 5686 -4172 6374 -3748
rect 6438 -4172 6458 -3748
rect 5686 -4200 6458 -4172
rect 6698 -3748 7470 -3720
rect 6698 -4172 7386 -3748
rect 7450 -4172 7470 -3748
rect 6698 -4200 7470 -4172
rect -7470 -4468 -6698 -4440
rect -7470 -4892 -6782 -4468
rect -6718 -4892 -6698 -4468
rect -7470 -4920 -6698 -4892
rect -6458 -4468 -5686 -4440
rect -6458 -4892 -5770 -4468
rect -5706 -4892 -5686 -4468
rect -6458 -4920 -5686 -4892
rect -5446 -4468 -4674 -4440
rect -5446 -4892 -4758 -4468
rect -4694 -4892 -4674 -4468
rect -5446 -4920 -4674 -4892
rect -4434 -4468 -3662 -4440
rect -4434 -4892 -3746 -4468
rect -3682 -4892 -3662 -4468
rect -4434 -4920 -3662 -4892
rect -3422 -4468 -2650 -4440
rect -3422 -4892 -2734 -4468
rect -2670 -4892 -2650 -4468
rect -3422 -4920 -2650 -4892
rect -2410 -4468 -1638 -4440
rect -2410 -4892 -1722 -4468
rect -1658 -4892 -1638 -4468
rect -2410 -4920 -1638 -4892
rect -1398 -4468 -626 -4440
rect -1398 -4892 -710 -4468
rect -646 -4892 -626 -4468
rect -1398 -4920 -626 -4892
rect -386 -4468 386 -4440
rect -386 -4892 302 -4468
rect 366 -4892 386 -4468
rect -386 -4920 386 -4892
rect 626 -4468 1398 -4440
rect 626 -4892 1314 -4468
rect 1378 -4892 1398 -4468
rect 626 -4920 1398 -4892
rect 1638 -4468 2410 -4440
rect 1638 -4892 2326 -4468
rect 2390 -4892 2410 -4468
rect 1638 -4920 2410 -4892
rect 2650 -4468 3422 -4440
rect 2650 -4892 3338 -4468
rect 3402 -4892 3422 -4468
rect 2650 -4920 3422 -4892
rect 3662 -4468 4434 -4440
rect 3662 -4892 4350 -4468
rect 4414 -4892 4434 -4468
rect 3662 -4920 4434 -4892
rect 4674 -4468 5446 -4440
rect 4674 -4892 5362 -4468
rect 5426 -4892 5446 -4468
rect 4674 -4920 5446 -4892
rect 5686 -4468 6458 -4440
rect 5686 -4892 6374 -4468
rect 6438 -4892 6458 -4468
rect 5686 -4920 6458 -4892
rect 6698 -4468 7470 -4440
rect 6698 -4892 7386 -4468
rect 7450 -4892 7470 -4468
rect 6698 -4920 7470 -4892
rect -7470 -5188 -6698 -5160
rect -7470 -5612 -6782 -5188
rect -6718 -5612 -6698 -5188
rect -7470 -5640 -6698 -5612
rect -6458 -5188 -5686 -5160
rect -6458 -5612 -5770 -5188
rect -5706 -5612 -5686 -5188
rect -6458 -5640 -5686 -5612
rect -5446 -5188 -4674 -5160
rect -5446 -5612 -4758 -5188
rect -4694 -5612 -4674 -5188
rect -5446 -5640 -4674 -5612
rect -4434 -5188 -3662 -5160
rect -4434 -5612 -3746 -5188
rect -3682 -5612 -3662 -5188
rect -4434 -5640 -3662 -5612
rect -3422 -5188 -2650 -5160
rect -3422 -5612 -2734 -5188
rect -2670 -5612 -2650 -5188
rect -3422 -5640 -2650 -5612
rect -2410 -5188 -1638 -5160
rect -2410 -5612 -1722 -5188
rect -1658 -5612 -1638 -5188
rect -2410 -5640 -1638 -5612
rect -1398 -5188 -626 -5160
rect -1398 -5612 -710 -5188
rect -646 -5612 -626 -5188
rect -1398 -5640 -626 -5612
rect -386 -5188 386 -5160
rect -386 -5612 302 -5188
rect 366 -5612 386 -5188
rect -386 -5640 386 -5612
rect 626 -5188 1398 -5160
rect 626 -5612 1314 -5188
rect 1378 -5612 1398 -5188
rect 626 -5640 1398 -5612
rect 1638 -5188 2410 -5160
rect 1638 -5612 2326 -5188
rect 2390 -5612 2410 -5188
rect 1638 -5640 2410 -5612
rect 2650 -5188 3422 -5160
rect 2650 -5612 3338 -5188
rect 3402 -5612 3422 -5188
rect 2650 -5640 3422 -5612
rect 3662 -5188 4434 -5160
rect 3662 -5612 4350 -5188
rect 4414 -5612 4434 -5188
rect 3662 -5640 4434 -5612
rect 4674 -5188 5446 -5160
rect 4674 -5612 5362 -5188
rect 5426 -5612 5446 -5188
rect 4674 -5640 5446 -5612
rect 5686 -5188 6458 -5160
rect 5686 -5612 6374 -5188
rect 6438 -5612 6458 -5188
rect 5686 -5640 6458 -5612
rect 6698 -5188 7470 -5160
rect 6698 -5612 7386 -5188
rect 7450 -5612 7470 -5188
rect 6698 -5640 7470 -5612
rect -7470 -5908 -6698 -5880
rect -7470 -6332 -6782 -5908
rect -6718 -6332 -6698 -5908
rect -7470 -6360 -6698 -6332
rect -6458 -5908 -5686 -5880
rect -6458 -6332 -5770 -5908
rect -5706 -6332 -5686 -5908
rect -6458 -6360 -5686 -6332
rect -5446 -5908 -4674 -5880
rect -5446 -6332 -4758 -5908
rect -4694 -6332 -4674 -5908
rect -5446 -6360 -4674 -6332
rect -4434 -5908 -3662 -5880
rect -4434 -6332 -3746 -5908
rect -3682 -6332 -3662 -5908
rect -4434 -6360 -3662 -6332
rect -3422 -5908 -2650 -5880
rect -3422 -6332 -2734 -5908
rect -2670 -6332 -2650 -5908
rect -3422 -6360 -2650 -6332
rect -2410 -5908 -1638 -5880
rect -2410 -6332 -1722 -5908
rect -1658 -6332 -1638 -5908
rect -2410 -6360 -1638 -6332
rect -1398 -5908 -626 -5880
rect -1398 -6332 -710 -5908
rect -646 -6332 -626 -5908
rect -1398 -6360 -626 -6332
rect -386 -5908 386 -5880
rect -386 -6332 302 -5908
rect 366 -6332 386 -5908
rect -386 -6360 386 -6332
rect 626 -5908 1398 -5880
rect 626 -6332 1314 -5908
rect 1378 -6332 1398 -5908
rect 626 -6360 1398 -6332
rect 1638 -5908 2410 -5880
rect 1638 -6332 2326 -5908
rect 2390 -6332 2410 -5908
rect 1638 -6360 2410 -6332
rect 2650 -5908 3422 -5880
rect 2650 -6332 3338 -5908
rect 3402 -6332 3422 -5908
rect 2650 -6360 3422 -6332
rect 3662 -5908 4434 -5880
rect 3662 -6332 4350 -5908
rect 4414 -6332 4434 -5908
rect 3662 -6360 4434 -6332
rect 4674 -5908 5446 -5880
rect 4674 -6332 5362 -5908
rect 5426 -6332 5446 -5908
rect 4674 -6360 5446 -6332
rect 5686 -5908 6458 -5880
rect 5686 -6332 6374 -5908
rect 6438 -6332 6458 -5908
rect 5686 -6360 6458 -6332
rect 6698 -5908 7470 -5880
rect 6698 -6332 7386 -5908
rect 7450 -6332 7470 -5908
rect 6698 -6360 7470 -6332
rect -7470 -6628 -6698 -6600
rect -7470 -7052 -6782 -6628
rect -6718 -7052 -6698 -6628
rect -7470 -7080 -6698 -7052
rect -6458 -6628 -5686 -6600
rect -6458 -7052 -5770 -6628
rect -5706 -7052 -5686 -6628
rect -6458 -7080 -5686 -7052
rect -5446 -6628 -4674 -6600
rect -5446 -7052 -4758 -6628
rect -4694 -7052 -4674 -6628
rect -5446 -7080 -4674 -7052
rect -4434 -6628 -3662 -6600
rect -4434 -7052 -3746 -6628
rect -3682 -7052 -3662 -6628
rect -4434 -7080 -3662 -7052
rect -3422 -6628 -2650 -6600
rect -3422 -7052 -2734 -6628
rect -2670 -7052 -2650 -6628
rect -3422 -7080 -2650 -7052
rect -2410 -6628 -1638 -6600
rect -2410 -7052 -1722 -6628
rect -1658 -7052 -1638 -6628
rect -2410 -7080 -1638 -7052
rect -1398 -6628 -626 -6600
rect -1398 -7052 -710 -6628
rect -646 -7052 -626 -6628
rect -1398 -7080 -626 -7052
rect -386 -6628 386 -6600
rect -386 -7052 302 -6628
rect 366 -7052 386 -6628
rect -386 -7080 386 -7052
rect 626 -6628 1398 -6600
rect 626 -7052 1314 -6628
rect 1378 -7052 1398 -6628
rect 626 -7080 1398 -7052
rect 1638 -6628 2410 -6600
rect 1638 -7052 2326 -6628
rect 2390 -7052 2410 -6628
rect 1638 -7080 2410 -7052
rect 2650 -6628 3422 -6600
rect 2650 -7052 3338 -6628
rect 3402 -7052 3422 -6628
rect 2650 -7080 3422 -7052
rect 3662 -6628 4434 -6600
rect 3662 -7052 4350 -6628
rect 4414 -7052 4434 -6628
rect 3662 -7080 4434 -7052
rect 4674 -6628 5446 -6600
rect 4674 -7052 5362 -6628
rect 5426 -7052 5446 -6628
rect 4674 -7080 5446 -7052
rect 5686 -6628 6458 -6600
rect 5686 -7052 6374 -6628
rect 6438 -7052 6458 -6628
rect 5686 -7080 6458 -7052
rect 6698 -6628 7470 -6600
rect 6698 -7052 7386 -6628
rect 7450 -7052 7470 -6628
rect 6698 -7080 7470 -7052
rect -7470 -7348 -6698 -7320
rect -7470 -7772 -6782 -7348
rect -6718 -7772 -6698 -7348
rect -7470 -7800 -6698 -7772
rect -6458 -7348 -5686 -7320
rect -6458 -7772 -5770 -7348
rect -5706 -7772 -5686 -7348
rect -6458 -7800 -5686 -7772
rect -5446 -7348 -4674 -7320
rect -5446 -7772 -4758 -7348
rect -4694 -7772 -4674 -7348
rect -5446 -7800 -4674 -7772
rect -4434 -7348 -3662 -7320
rect -4434 -7772 -3746 -7348
rect -3682 -7772 -3662 -7348
rect -4434 -7800 -3662 -7772
rect -3422 -7348 -2650 -7320
rect -3422 -7772 -2734 -7348
rect -2670 -7772 -2650 -7348
rect -3422 -7800 -2650 -7772
rect -2410 -7348 -1638 -7320
rect -2410 -7772 -1722 -7348
rect -1658 -7772 -1638 -7348
rect -2410 -7800 -1638 -7772
rect -1398 -7348 -626 -7320
rect -1398 -7772 -710 -7348
rect -646 -7772 -626 -7348
rect -1398 -7800 -626 -7772
rect -386 -7348 386 -7320
rect -386 -7772 302 -7348
rect 366 -7772 386 -7348
rect -386 -7800 386 -7772
rect 626 -7348 1398 -7320
rect 626 -7772 1314 -7348
rect 1378 -7772 1398 -7348
rect 626 -7800 1398 -7772
rect 1638 -7348 2410 -7320
rect 1638 -7772 2326 -7348
rect 2390 -7772 2410 -7348
rect 1638 -7800 2410 -7772
rect 2650 -7348 3422 -7320
rect 2650 -7772 3338 -7348
rect 3402 -7772 3422 -7348
rect 2650 -7800 3422 -7772
rect 3662 -7348 4434 -7320
rect 3662 -7772 4350 -7348
rect 4414 -7772 4434 -7348
rect 3662 -7800 4434 -7772
rect 4674 -7348 5446 -7320
rect 4674 -7772 5362 -7348
rect 5426 -7772 5446 -7348
rect 4674 -7800 5446 -7772
rect 5686 -7348 6458 -7320
rect 5686 -7772 6374 -7348
rect 6438 -7772 6458 -7348
rect 5686 -7800 6458 -7772
rect 6698 -7348 7470 -7320
rect 6698 -7772 7386 -7348
rect 7450 -7772 7470 -7348
rect 6698 -7800 7470 -7772
rect -7470 -8068 -6698 -8040
rect -7470 -8492 -6782 -8068
rect -6718 -8492 -6698 -8068
rect -7470 -8520 -6698 -8492
rect -6458 -8068 -5686 -8040
rect -6458 -8492 -5770 -8068
rect -5706 -8492 -5686 -8068
rect -6458 -8520 -5686 -8492
rect -5446 -8068 -4674 -8040
rect -5446 -8492 -4758 -8068
rect -4694 -8492 -4674 -8068
rect -5446 -8520 -4674 -8492
rect -4434 -8068 -3662 -8040
rect -4434 -8492 -3746 -8068
rect -3682 -8492 -3662 -8068
rect -4434 -8520 -3662 -8492
rect -3422 -8068 -2650 -8040
rect -3422 -8492 -2734 -8068
rect -2670 -8492 -2650 -8068
rect -3422 -8520 -2650 -8492
rect -2410 -8068 -1638 -8040
rect -2410 -8492 -1722 -8068
rect -1658 -8492 -1638 -8068
rect -2410 -8520 -1638 -8492
rect -1398 -8068 -626 -8040
rect -1398 -8492 -710 -8068
rect -646 -8492 -626 -8068
rect -1398 -8520 -626 -8492
rect -386 -8068 386 -8040
rect -386 -8492 302 -8068
rect 366 -8492 386 -8068
rect -386 -8520 386 -8492
rect 626 -8068 1398 -8040
rect 626 -8492 1314 -8068
rect 1378 -8492 1398 -8068
rect 626 -8520 1398 -8492
rect 1638 -8068 2410 -8040
rect 1638 -8492 2326 -8068
rect 2390 -8492 2410 -8068
rect 1638 -8520 2410 -8492
rect 2650 -8068 3422 -8040
rect 2650 -8492 3338 -8068
rect 3402 -8492 3422 -8068
rect 2650 -8520 3422 -8492
rect 3662 -8068 4434 -8040
rect 3662 -8492 4350 -8068
rect 4414 -8492 4434 -8068
rect 3662 -8520 4434 -8492
rect 4674 -8068 5446 -8040
rect 4674 -8492 5362 -8068
rect 5426 -8492 5446 -8068
rect 4674 -8520 5446 -8492
rect 5686 -8068 6458 -8040
rect 5686 -8492 6374 -8068
rect 6438 -8492 6458 -8068
rect 5686 -8520 6458 -8492
rect 6698 -8068 7470 -8040
rect 6698 -8492 7386 -8068
rect 7450 -8492 7470 -8068
rect 6698 -8520 7470 -8492
rect -7470 -8788 -6698 -8760
rect -7470 -9212 -6782 -8788
rect -6718 -9212 -6698 -8788
rect -7470 -9240 -6698 -9212
rect -6458 -8788 -5686 -8760
rect -6458 -9212 -5770 -8788
rect -5706 -9212 -5686 -8788
rect -6458 -9240 -5686 -9212
rect -5446 -8788 -4674 -8760
rect -5446 -9212 -4758 -8788
rect -4694 -9212 -4674 -8788
rect -5446 -9240 -4674 -9212
rect -4434 -8788 -3662 -8760
rect -4434 -9212 -3746 -8788
rect -3682 -9212 -3662 -8788
rect -4434 -9240 -3662 -9212
rect -3422 -8788 -2650 -8760
rect -3422 -9212 -2734 -8788
rect -2670 -9212 -2650 -8788
rect -3422 -9240 -2650 -9212
rect -2410 -8788 -1638 -8760
rect -2410 -9212 -1722 -8788
rect -1658 -9212 -1638 -8788
rect -2410 -9240 -1638 -9212
rect -1398 -8788 -626 -8760
rect -1398 -9212 -710 -8788
rect -646 -9212 -626 -8788
rect -1398 -9240 -626 -9212
rect -386 -8788 386 -8760
rect -386 -9212 302 -8788
rect 366 -9212 386 -8788
rect -386 -9240 386 -9212
rect 626 -8788 1398 -8760
rect 626 -9212 1314 -8788
rect 1378 -9212 1398 -8788
rect 626 -9240 1398 -9212
rect 1638 -8788 2410 -8760
rect 1638 -9212 2326 -8788
rect 2390 -9212 2410 -8788
rect 1638 -9240 2410 -9212
rect 2650 -8788 3422 -8760
rect 2650 -9212 3338 -8788
rect 3402 -9212 3422 -8788
rect 2650 -9240 3422 -9212
rect 3662 -8788 4434 -8760
rect 3662 -9212 4350 -8788
rect 4414 -9212 4434 -8788
rect 3662 -9240 4434 -9212
rect 4674 -8788 5446 -8760
rect 4674 -9212 5362 -8788
rect 5426 -9212 5446 -8788
rect 4674 -9240 5446 -9212
rect 5686 -8788 6458 -8760
rect 5686 -9212 6374 -8788
rect 6438 -9212 6458 -8788
rect 5686 -9240 6458 -9212
rect 6698 -8788 7470 -8760
rect 6698 -9212 7386 -8788
rect 7450 -9212 7470 -8788
rect 6698 -9240 7470 -9212
rect -7470 -9508 -6698 -9480
rect -7470 -9932 -6782 -9508
rect -6718 -9932 -6698 -9508
rect -7470 -9960 -6698 -9932
rect -6458 -9508 -5686 -9480
rect -6458 -9932 -5770 -9508
rect -5706 -9932 -5686 -9508
rect -6458 -9960 -5686 -9932
rect -5446 -9508 -4674 -9480
rect -5446 -9932 -4758 -9508
rect -4694 -9932 -4674 -9508
rect -5446 -9960 -4674 -9932
rect -4434 -9508 -3662 -9480
rect -4434 -9932 -3746 -9508
rect -3682 -9932 -3662 -9508
rect -4434 -9960 -3662 -9932
rect -3422 -9508 -2650 -9480
rect -3422 -9932 -2734 -9508
rect -2670 -9932 -2650 -9508
rect -3422 -9960 -2650 -9932
rect -2410 -9508 -1638 -9480
rect -2410 -9932 -1722 -9508
rect -1658 -9932 -1638 -9508
rect -2410 -9960 -1638 -9932
rect -1398 -9508 -626 -9480
rect -1398 -9932 -710 -9508
rect -646 -9932 -626 -9508
rect -1398 -9960 -626 -9932
rect -386 -9508 386 -9480
rect -386 -9932 302 -9508
rect 366 -9932 386 -9508
rect -386 -9960 386 -9932
rect 626 -9508 1398 -9480
rect 626 -9932 1314 -9508
rect 1378 -9932 1398 -9508
rect 626 -9960 1398 -9932
rect 1638 -9508 2410 -9480
rect 1638 -9932 2326 -9508
rect 2390 -9932 2410 -9508
rect 1638 -9960 2410 -9932
rect 2650 -9508 3422 -9480
rect 2650 -9932 3338 -9508
rect 3402 -9932 3422 -9508
rect 2650 -9960 3422 -9932
rect 3662 -9508 4434 -9480
rect 3662 -9932 4350 -9508
rect 4414 -9932 4434 -9508
rect 3662 -9960 4434 -9932
rect 4674 -9508 5446 -9480
rect 4674 -9932 5362 -9508
rect 5426 -9932 5446 -9508
rect 4674 -9960 5446 -9932
rect 5686 -9508 6458 -9480
rect 5686 -9932 6374 -9508
rect 6438 -9932 6458 -9508
rect 5686 -9960 6458 -9932
rect 6698 -9508 7470 -9480
rect 6698 -9932 7386 -9508
rect 7450 -9932 7470 -9508
rect 6698 -9960 7470 -9932
rect -7470 -10228 -6698 -10200
rect -7470 -10652 -6782 -10228
rect -6718 -10652 -6698 -10228
rect -7470 -10680 -6698 -10652
rect -6458 -10228 -5686 -10200
rect -6458 -10652 -5770 -10228
rect -5706 -10652 -5686 -10228
rect -6458 -10680 -5686 -10652
rect -5446 -10228 -4674 -10200
rect -5446 -10652 -4758 -10228
rect -4694 -10652 -4674 -10228
rect -5446 -10680 -4674 -10652
rect -4434 -10228 -3662 -10200
rect -4434 -10652 -3746 -10228
rect -3682 -10652 -3662 -10228
rect -4434 -10680 -3662 -10652
rect -3422 -10228 -2650 -10200
rect -3422 -10652 -2734 -10228
rect -2670 -10652 -2650 -10228
rect -3422 -10680 -2650 -10652
rect -2410 -10228 -1638 -10200
rect -2410 -10652 -1722 -10228
rect -1658 -10652 -1638 -10228
rect -2410 -10680 -1638 -10652
rect -1398 -10228 -626 -10200
rect -1398 -10652 -710 -10228
rect -646 -10652 -626 -10228
rect -1398 -10680 -626 -10652
rect -386 -10228 386 -10200
rect -386 -10652 302 -10228
rect 366 -10652 386 -10228
rect -386 -10680 386 -10652
rect 626 -10228 1398 -10200
rect 626 -10652 1314 -10228
rect 1378 -10652 1398 -10228
rect 626 -10680 1398 -10652
rect 1638 -10228 2410 -10200
rect 1638 -10652 2326 -10228
rect 2390 -10652 2410 -10228
rect 1638 -10680 2410 -10652
rect 2650 -10228 3422 -10200
rect 2650 -10652 3338 -10228
rect 3402 -10652 3422 -10228
rect 2650 -10680 3422 -10652
rect 3662 -10228 4434 -10200
rect 3662 -10652 4350 -10228
rect 4414 -10652 4434 -10228
rect 3662 -10680 4434 -10652
rect 4674 -10228 5446 -10200
rect 4674 -10652 5362 -10228
rect 5426 -10652 5446 -10228
rect 4674 -10680 5446 -10652
rect 5686 -10228 6458 -10200
rect 5686 -10652 6374 -10228
rect 6438 -10652 6458 -10228
rect 5686 -10680 6458 -10652
rect 6698 -10228 7470 -10200
rect 6698 -10652 7386 -10228
rect 7450 -10652 7470 -10228
rect 6698 -10680 7470 -10652
rect -7470 -10948 -6698 -10920
rect -7470 -11372 -6782 -10948
rect -6718 -11372 -6698 -10948
rect -7470 -11400 -6698 -11372
rect -6458 -10948 -5686 -10920
rect -6458 -11372 -5770 -10948
rect -5706 -11372 -5686 -10948
rect -6458 -11400 -5686 -11372
rect -5446 -10948 -4674 -10920
rect -5446 -11372 -4758 -10948
rect -4694 -11372 -4674 -10948
rect -5446 -11400 -4674 -11372
rect -4434 -10948 -3662 -10920
rect -4434 -11372 -3746 -10948
rect -3682 -11372 -3662 -10948
rect -4434 -11400 -3662 -11372
rect -3422 -10948 -2650 -10920
rect -3422 -11372 -2734 -10948
rect -2670 -11372 -2650 -10948
rect -3422 -11400 -2650 -11372
rect -2410 -10948 -1638 -10920
rect -2410 -11372 -1722 -10948
rect -1658 -11372 -1638 -10948
rect -2410 -11400 -1638 -11372
rect -1398 -10948 -626 -10920
rect -1398 -11372 -710 -10948
rect -646 -11372 -626 -10948
rect -1398 -11400 -626 -11372
rect -386 -10948 386 -10920
rect -386 -11372 302 -10948
rect 366 -11372 386 -10948
rect -386 -11400 386 -11372
rect 626 -10948 1398 -10920
rect 626 -11372 1314 -10948
rect 1378 -11372 1398 -10948
rect 626 -11400 1398 -11372
rect 1638 -10948 2410 -10920
rect 1638 -11372 2326 -10948
rect 2390 -11372 2410 -10948
rect 1638 -11400 2410 -11372
rect 2650 -10948 3422 -10920
rect 2650 -11372 3338 -10948
rect 3402 -11372 3422 -10948
rect 2650 -11400 3422 -11372
rect 3662 -10948 4434 -10920
rect 3662 -11372 4350 -10948
rect 4414 -11372 4434 -10948
rect 3662 -11400 4434 -11372
rect 4674 -10948 5446 -10920
rect 4674 -11372 5362 -10948
rect 5426 -11372 5446 -10948
rect 4674 -11400 5446 -11372
rect 5686 -10948 6458 -10920
rect 5686 -11372 6374 -10948
rect 6438 -11372 6458 -10948
rect 5686 -11400 6458 -11372
rect 6698 -10948 7470 -10920
rect 6698 -11372 7386 -10948
rect 7450 -11372 7470 -10948
rect 6698 -11400 7470 -11372
<< via3 >>
rect -6782 10948 -6718 11372
rect -5770 10948 -5706 11372
rect -4758 10948 -4694 11372
rect -3746 10948 -3682 11372
rect -2734 10948 -2670 11372
rect -1722 10948 -1658 11372
rect -710 10948 -646 11372
rect 302 10948 366 11372
rect 1314 10948 1378 11372
rect 2326 10948 2390 11372
rect 3338 10948 3402 11372
rect 4350 10948 4414 11372
rect 5362 10948 5426 11372
rect 6374 10948 6438 11372
rect 7386 10948 7450 11372
rect -6782 10228 -6718 10652
rect -5770 10228 -5706 10652
rect -4758 10228 -4694 10652
rect -3746 10228 -3682 10652
rect -2734 10228 -2670 10652
rect -1722 10228 -1658 10652
rect -710 10228 -646 10652
rect 302 10228 366 10652
rect 1314 10228 1378 10652
rect 2326 10228 2390 10652
rect 3338 10228 3402 10652
rect 4350 10228 4414 10652
rect 5362 10228 5426 10652
rect 6374 10228 6438 10652
rect 7386 10228 7450 10652
rect -6782 9508 -6718 9932
rect -5770 9508 -5706 9932
rect -4758 9508 -4694 9932
rect -3746 9508 -3682 9932
rect -2734 9508 -2670 9932
rect -1722 9508 -1658 9932
rect -710 9508 -646 9932
rect 302 9508 366 9932
rect 1314 9508 1378 9932
rect 2326 9508 2390 9932
rect 3338 9508 3402 9932
rect 4350 9508 4414 9932
rect 5362 9508 5426 9932
rect 6374 9508 6438 9932
rect 7386 9508 7450 9932
rect -6782 8788 -6718 9212
rect -5770 8788 -5706 9212
rect -4758 8788 -4694 9212
rect -3746 8788 -3682 9212
rect -2734 8788 -2670 9212
rect -1722 8788 -1658 9212
rect -710 8788 -646 9212
rect 302 8788 366 9212
rect 1314 8788 1378 9212
rect 2326 8788 2390 9212
rect 3338 8788 3402 9212
rect 4350 8788 4414 9212
rect 5362 8788 5426 9212
rect 6374 8788 6438 9212
rect 7386 8788 7450 9212
rect -6782 8068 -6718 8492
rect -5770 8068 -5706 8492
rect -4758 8068 -4694 8492
rect -3746 8068 -3682 8492
rect -2734 8068 -2670 8492
rect -1722 8068 -1658 8492
rect -710 8068 -646 8492
rect 302 8068 366 8492
rect 1314 8068 1378 8492
rect 2326 8068 2390 8492
rect 3338 8068 3402 8492
rect 4350 8068 4414 8492
rect 5362 8068 5426 8492
rect 6374 8068 6438 8492
rect 7386 8068 7450 8492
rect -6782 7348 -6718 7772
rect -5770 7348 -5706 7772
rect -4758 7348 -4694 7772
rect -3746 7348 -3682 7772
rect -2734 7348 -2670 7772
rect -1722 7348 -1658 7772
rect -710 7348 -646 7772
rect 302 7348 366 7772
rect 1314 7348 1378 7772
rect 2326 7348 2390 7772
rect 3338 7348 3402 7772
rect 4350 7348 4414 7772
rect 5362 7348 5426 7772
rect 6374 7348 6438 7772
rect 7386 7348 7450 7772
rect -6782 6628 -6718 7052
rect -5770 6628 -5706 7052
rect -4758 6628 -4694 7052
rect -3746 6628 -3682 7052
rect -2734 6628 -2670 7052
rect -1722 6628 -1658 7052
rect -710 6628 -646 7052
rect 302 6628 366 7052
rect 1314 6628 1378 7052
rect 2326 6628 2390 7052
rect 3338 6628 3402 7052
rect 4350 6628 4414 7052
rect 5362 6628 5426 7052
rect 6374 6628 6438 7052
rect 7386 6628 7450 7052
rect -6782 5908 -6718 6332
rect -5770 5908 -5706 6332
rect -4758 5908 -4694 6332
rect -3746 5908 -3682 6332
rect -2734 5908 -2670 6332
rect -1722 5908 -1658 6332
rect -710 5908 -646 6332
rect 302 5908 366 6332
rect 1314 5908 1378 6332
rect 2326 5908 2390 6332
rect 3338 5908 3402 6332
rect 4350 5908 4414 6332
rect 5362 5908 5426 6332
rect 6374 5908 6438 6332
rect 7386 5908 7450 6332
rect -6782 5188 -6718 5612
rect -5770 5188 -5706 5612
rect -4758 5188 -4694 5612
rect -3746 5188 -3682 5612
rect -2734 5188 -2670 5612
rect -1722 5188 -1658 5612
rect -710 5188 -646 5612
rect 302 5188 366 5612
rect 1314 5188 1378 5612
rect 2326 5188 2390 5612
rect 3338 5188 3402 5612
rect 4350 5188 4414 5612
rect 5362 5188 5426 5612
rect 6374 5188 6438 5612
rect 7386 5188 7450 5612
rect -6782 4468 -6718 4892
rect -5770 4468 -5706 4892
rect -4758 4468 -4694 4892
rect -3746 4468 -3682 4892
rect -2734 4468 -2670 4892
rect -1722 4468 -1658 4892
rect -710 4468 -646 4892
rect 302 4468 366 4892
rect 1314 4468 1378 4892
rect 2326 4468 2390 4892
rect 3338 4468 3402 4892
rect 4350 4468 4414 4892
rect 5362 4468 5426 4892
rect 6374 4468 6438 4892
rect 7386 4468 7450 4892
rect -6782 3748 -6718 4172
rect -5770 3748 -5706 4172
rect -4758 3748 -4694 4172
rect -3746 3748 -3682 4172
rect -2734 3748 -2670 4172
rect -1722 3748 -1658 4172
rect -710 3748 -646 4172
rect 302 3748 366 4172
rect 1314 3748 1378 4172
rect 2326 3748 2390 4172
rect 3338 3748 3402 4172
rect 4350 3748 4414 4172
rect 5362 3748 5426 4172
rect 6374 3748 6438 4172
rect 7386 3748 7450 4172
rect -6782 3028 -6718 3452
rect -5770 3028 -5706 3452
rect -4758 3028 -4694 3452
rect -3746 3028 -3682 3452
rect -2734 3028 -2670 3452
rect -1722 3028 -1658 3452
rect -710 3028 -646 3452
rect 302 3028 366 3452
rect 1314 3028 1378 3452
rect 2326 3028 2390 3452
rect 3338 3028 3402 3452
rect 4350 3028 4414 3452
rect 5362 3028 5426 3452
rect 6374 3028 6438 3452
rect 7386 3028 7450 3452
rect -6782 2308 -6718 2732
rect -5770 2308 -5706 2732
rect -4758 2308 -4694 2732
rect -3746 2308 -3682 2732
rect -2734 2308 -2670 2732
rect -1722 2308 -1658 2732
rect -710 2308 -646 2732
rect 302 2308 366 2732
rect 1314 2308 1378 2732
rect 2326 2308 2390 2732
rect 3338 2308 3402 2732
rect 4350 2308 4414 2732
rect 5362 2308 5426 2732
rect 6374 2308 6438 2732
rect 7386 2308 7450 2732
rect -6782 1588 -6718 2012
rect -5770 1588 -5706 2012
rect -4758 1588 -4694 2012
rect -3746 1588 -3682 2012
rect -2734 1588 -2670 2012
rect -1722 1588 -1658 2012
rect -710 1588 -646 2012
rect 302 1588 366 2012
rect 1314 1588 1378 2012
rect 2326 1588 2390 2012
rect 3338 1588 3402 2012
rect 4350 1588 4414 2012
rect 5362 1588 5426 2012
rect 6374 1588 6438 2012
rect 7386 1588 7450 2012
rect -6782 868 -6718 1292
rect -5770 868 -5706 1292
rect -4758 868 -4694 1292
rect -3746 868 -3682 1292
rect -2734 868 -2670 1292
rect -1722 868 -1658 1292
rect -710 868 -646 1292
rect 302 868 366 1292
rect 1314 868 1378 1292
rect 2326 868 2390 1292
rect 3338 868 3402 1292
rect 4350 868 4414 1292
rect 5362 868 5426 1292
rect 6374 868 6438 1292
rect 7386 868 7450 1292
rect -6782 148 -6718 572
rect -5770 148 -5706 572
rect -4758 148 -4694 572
rect -3746 148 -3682 572
rect -2734 148 -2670 572
rect -1722 148 -1658 572
rect -710 148 -646 572
rect 302 148 366 572
rect 1314 148 1378 572
rect 2326 148 2390 572
rect 3338 148 3402 572
rect 4350 148 4414 572
rect 5362 148 5426 572
rect 6374 148 6438 572
rect 7386 148 7450 572
rect -6782 -572 -6718 -148
rect -5770 -572 -5706 -148
rect -4758 -572 -4694 -148
rect -3746 -572 -3682 -148
rect -2734 -572 -2670 -148
rect -1722 -572 -1658 -148
rect -710 -572 -646 -148
rect 302 -572 366 -148
rect 1314 -572 1378 -148
rect 2326 -572 2390 -148
rect 3338 -572 3402 -148
rect 4350 -572 4414 -148
rect 5362 -572 5426 -148
rect 6374 -572 6438 -148
rect 7386 -572 7450 -148
rect -6782 -1292 -6718 -868
rect -5770 -1292 -5706 -868
rect -4758 -1292 -4694 -868
rect -3746 -1292 -3682 -868
rect -2734 -1292 -2670 -868
rect -1722 -1292 -1658 -868
rect -710 -1292 -646 -868
rect 302 -1292 366 -868
rect 1314 -1292 1378 -868
rect 2326 -1292 2390 -868
rect 3338 -1292 3402 -868
rect 4350 -1292 4414 -868
rect 5362 -1292 5426 -868
rect 6374 -1292 6438 -868
rect 7386 -1292 7450 -868
rect -6782 -2012 -6718 -1588
rect -5770 -2012 -5706 -1588
rect -4758 -2012 -4694 -1588
rect -3746 -2012 -3682 -1588
rect -2734 -2012 -2670 -1588
rect -1722 -2012 -1658 -1588
rect -710 -2012 -646 -1588
rect 302 -2012 366 -1588
rect 1314 -2012 1378 -1588
rect 2326 -2012 2390 -1588
rect 3338 -2012 3402 -1588
rect 4350 -2012 4414 -1588
rect 5362 -2012 5426 -1588
rect 6374 -2012 6438 -1588
rect 7386 -2012 7450 -1588
rect -6782 -2732 -6718 -2308
rect -5770 -2732 -5706 -2308
rect -4758 -2732 -4694 -2308
rect -3746 -2732 -3682 -2308
rect -2734 -2732 -2670 -2308
rect -1722 -2732 -1658 -2308
rect -710 -2732 -646 -2308
rect 302 -2732 366 -2308
rect 1314 -2732 1378 -2308
rect 2326 -2732 2390 -2308
rect 3338 -2732 3402 -2308
rect 4350 -2732 4414 -2308
rect 5362 -2732 5426 -2308
rect 6374 -2732 6438 -2308
rect 7386 -2732 7450 -2308
rect -6782 -3452 -6718 -3028
rect -5770 -3452 -5706 -3028
rect -4758 -3452 -4694 -3028
rect -3746 -3452 -3682 -3028
rect -2734 -3452 -2670 -3028
rect -1722 -3452 -1658 -3028
rect -710 -3452 -646 -3028
rect 302 -3452 366 -3028
rect 1314 -3452 1378 -3028
rect 2326 -3452 2390 -3028
rect 3338 -3452 3402 -3028
rect 4350 -3452 4414 -3028
rect 5362 -3452 5426 -3028
rect 6374 -3452 6438 -3028
rect 7386 -3452 7450 -3028
rect -6782 -4172 -6718 -3748
rect -5770 -4172 -5706 -3748
rect -4758 -4172 -4694 -3748
rect -3746 -4172 -3682 -3748
rect -2734 -4172 -2670 -3748
rect -1722 -4172 -1658 -3748
rect -710 -4172 -646 -3748
rect 302 -4172 366 -3748
rect 1314 -4172 1378 -3748
rect 2326 -4172 2390 -3748
rect 3338 -4172 3402 -3748
rect 4350 -4172 4414 -3748
rect 5362 -4172 5426 -3748
rect 6374 -4172 6438 -3748
rect 7386 -4172 7450 -3748
rect -6782 -4892 -6718 -4468
rect -5770 -4892 -5706 -4468
rect -4758 -4892 -4694 -4468
rect -3746 -4892 -3682 -4468
rect -2734 -4892 -2670 -4468
rect -1722 -4892 -1658 -4468
rect -710 -4892 -646 -4468
rect 302 -4892 366 -4468
rect 1314 -4892 1378 -4468
rect 2326 -4892 2390 -4468
rect 3338 -4892 3402 -4468
rect 4350 -4892 4414 -4468
rect 5362 -4892 5426 -4468
rect 6374 -4892 6438 -4468
rect 7386 -4892 7450 -4468
rect -6782 -5612 -6718 -5188
rect -5770 -5612 -5706 -5188
rect -4758 -5612 -4694 -5188
rect -3746 -5612 -3682 -5188
rect -2734 -5612 -2670 -5188
rect -1722 -5612 -1658 -5188
rect -710 -5612 -646 -5188
rect 302 -5612 366 -5188
rect 1314 -5612 1378 -5188
rect 2326 -5612 2390 -5188
rect 3338 -5612 3402 -5188
rect 4350 -5612 4414 -5188
rect 5362 -5612 5426 -5188
rect 6374 -5612 6438 -5188
rect 7386 -5612 7450 -5188
rect -6782 -6332 -6718 -5908
rect -5770 -6332 -5706 -5908
rect -4758 -6332 -4694 -5908
rect -3746 -6332 -3682 -5908
rect -2734 -6332 -2670 -5908
rect -1722 -6332 -1658 -5908
rect -710 -6332 -646 -5908
rect 302 -6332 366 -5908
rect 1314 -6332 1378 -5908
rect 2326 -6332 2390 -5908
rect 3338 -6332 3402 -5908
rect 4350 -6332 4414 -5908
rect 5362 -6332 5426 -5908
rect 6374 -6332 6438 -5908
rect 7386 -6332 7450 -5908
rect -6782 -7052 -6718 -6628
rect -5770 -7052 -5706 -6628
rect -4758 -7052 -4694 -6628
rect -3746 -7052 -3682 -6628
rect -2734 -7052 -2670 -6628
rect -1722 -7052 -1658 -6628
rect -710 -7052 -646 -6628
rect 302 -7052 366 -6628
rect 1314 -7052 1378 -6628
rect 2326 -7052 2390 -6628
rect 3338 -7052 3402 -6628
rect 4350 -7052 4414 -6628
rect 5362 -7052 5426 -6628
rect 6374 -7052 6438 -6628
rect 7386 -7052 7450 -6628
rect -6782 -7772 -6718 -7348
rect -5770 -7772 -5706 -7348
rect -4758 -7772 -4694 -7348
rect -3746 -7772 -3682 -7348
rect -2734 -7772 -2670 -7348
rect -1722 -7772 -1658 -7348
rect -710 -7772 -646 -7348
rect 302 -7772 366 -7348
rect 1314 -7772 1378 -7348
rect 2326 -7772 2390 -7348
rect 3338 -7772 3402 -7348
rect 4350 -7772 4414 -7348
rect 5362 -7772 5426 -7348
rect 6374 -7772 6438 -7348
rect 7386 -7772 7450 -7348
rect -6782 -8492 -6718 -8068
rect -5770 -8492 -5706 -8068
rect -4758 -8492 -4694 -8068
rect -3746 -8492 -3682 -8068
rect -2734 -8492 -2670 -8068
rect -1722 -8492 -1658 -8068
rect -710 -8492 -646 -8068
rect 302 -8492 366 -8068
rect 1314 -8492 1378 -8068
rect 2326 -8492 2390 -8068
rect 3338 -8492 3402 -8068
rect 4350 -8492 4414 -8068
rect 5362 -8492 5426 -8068
rect 6374 -8492 6438 -8068
rect 7386 -8492 7450 -8068
rect -6782 -9212 -6718 -8788
rect -5770 -9212 -5706 -8788
rect -4758 -9212 -4694 -8788
rect -3746 -9212 -3682 -8788
rect -2734 -9212 -2670 -8788
rect -1722 -9212 -1658 -8788
rect -710 -9212 -646 -8788
rect 302 -9212 366 -8788
rect 1314 -9212 1378 -8788
rect 2326 -9212 2390 -8788
rect 3338 -9212 3402 -8788
rect 4350 -9212 4414 -8788
rect 5362 -9212 5426 -8788
rect 6374 -9212 6438 -8788
rect 7386 -9212 7450 -8788
rect -6782 -9932 -6718 -9508
rect -5770 -9932 -5706 -9508
rect -4758 -9932 -4694 -9508
rect -3746 -9932 -3682 -9508
rect -2734 -9932 -2670 -9508
rect -1722 -9932 -1658 -9508
rect -710 -9932 -646 -9508
rect 302 -9932 366 -9508
rect 1314 -9932 1378 -9508
rect 2326 -9932 2390 -9508
rect 3338 -9932 3402 -9508
rect 4350 -9932 4414 -9508
rect 5362 -9932 5426 -9508
rect 6374 -9932 6438 -9508
rect 7386 -9932 7450 -9508
rect -6782 -10652 -6718 -10228
rect -5770 -10652 -5706 -10228
rect -4758 -10652 -4694 -10228
rect -3746 -10652 -3682 -10228
rect -2734 -10652 -2670 -10228
rect -1722 -10652 -1658 -10228
rect -710 -10652 -646 -10228
rect 302 -10652 366 -10228
rect 1314 -10652 1378 -10228
rect 2326 -10652 2390 -10228
rect 3338 -10652 3402 -10228
rect 4350 -10652 4414 -10228
rect 5362 -10652 5426 -10228
rect 6374 -10652 6438 -10228
rect 7386 -10652 7450 -10228
rect -6782 -11372 -6718 -10948
rect -5770 -11372 -5706 -10948
rect -4758 -11372 -4694 -10948
rect -3746 -11372 -3682 -10948
rect -2734 -11372 -2670 -10948
rect -1722 -11372 -1658 -10948
rect -710 -11372 -646 -10948
rect 302 -11372 366 -10948
rect 1314 -11372 1378 -10948
rect 2326 -11372 2390 -10948
rect 3338 -11372 3402 -10948
rect 4350 -11372 4414 -10948
rect 5362 -11372 5426 -10948
rect 6374 -11372 6438 -10948
rect 7386 -11372 7450 -10948
<< mimcap >>
rect -7430 11320 -7030 11360
rect -7430 11000 -7390 11320
rect -7070 11000 -7030 11320
rect -7430 10960 -7030 11000
rect -6418 11320 -6018 11360
rect -6418 11000 -6378 11320
rect -6058 11000 -6018 11320
rect -6418 10960 -6018 11000
rect -5406 11320 -5006 11360
rect -5406 11000 -5366 11320
rect -5046 11000 -5006 11320
rect -5406 10960 -5006 11000
rect -4394 11320 -3994 11360
rect -4394 11000 -4354 11320
rect -4034 11000 -3994 11320
rect -4394 10960 -3994 11000
rect -3382 11320 -2982 11360
rect -3382 11000 -3342 11320
rect -3022 11000 -2982 11320
rect -3382 10960 -2982 11000
rect -2370 11320 -1970 11360
rect -2370 11000 -2330 11320
rect -2010 11000 -1970 11320
rect -2370 10960 -1970 11000
rect -1358 11320 -958 11360
rect -1358 11000 -1318 11320
rect -998 11000 -958 11320
rect -1358 10960 -958 11000
rect -346 11320 54 11360
rect -346 11000 -306 11320
rect 14 11000 54 11320
rect -346 10960 54 11000
rect 666 11320 1066 11360
rect 666 11000 706 11320
rect 1026 11000 1066 11320
rect 666 10960 1066 11000
rect 1678 11320 2078 11360
rect 1678 11000 1718 11320
rect 2038 11000 2078 11320
rect 1678 10960 2078 11000
rect 2690 11320 3090 11360
rect 2690 11000 2730 11320
rect 3050 11000 3090 11320
rect 2690 10960 3090 11000
rect 3702 11320 4102 11360
rect 3702 11000 3742 11320
rect 4062 11000 4102 11320
rect 3702 10960 4102 11000
rect 4714 11320 5114 11360
rect 4714 11000 4754 11320
rect 5074 11000 5114 11320
rect 4714 10960 5114 11000
rect 5726 11320 6126 11360
rect 5726 11000 5766 11320
rect 6086 11000 6126 11320
rect 5726 10960 6126 11000
rect 6738 11320 7138 11360
rect 6738 11000 6778 11320
rect 7098 11000 7138 11320
rect 6738 10960 7138 11000
rect -7430 10600 -7030 10640
rect -7430 10280 -7390 10600
rect -7070 10280 -7030 10600
rect -7430 10240 -7030 10280
rect -6418 10600 -6018 10640
rect -6418 10280 -6378 10600
rect -6058 10280 -6018 10600
rect -6418 10240 -6018 10280
rect -5406 10600 -5006 10640
rect -5406 10280 -5366 10600
rect -5046 10280 -5006 10600
rect -5406 10240 -5006 10280
rect -4394 10600 -3994 10640
rect -4394 10280 -4354 10600
rect -4034 10280 -3994 10600
rect -4394 10240 -3994 10280
rect -3382 10600 -2982 10640
rect -3382 10280 -3342 10600
rect -3022 10280 -2982 10600
rect -3382 10240 -2982 10280
rect -2370 10600 -1970 10640
rect -2370 10280 -2330 10600
rect -2010 10280 -1970 10600
rect -2370 10240 -1970 10280
rect -1358 10600 -958 10640
rect -1358 10280 -1318 10600
rect -998 10280 -958 10600
rect -1358 10240 -958 10280
rect -346 10600 54 10640
rect -346 10280 -306 10600
rect 14 10280 54 10600
rect -346 10240 54 10280
rect 666 10600 1066 10640
rect 666 10280 706 10600
rect 1026 10280 1066 10600
rect 666 10240 1066 10280
rect 1678 10600 2078 10640
rect 1678 10280 1718 10600
rect 2038 10280 2078 10600
rect 1678 10240 2078 10280
rect 2690 10600 3090 10640
rect 2690 10280 2730 10600
rect 3050 10280 3090 10600
rect 2690 10240 3090 10280
rect 3702 10600 4102 10640
rect 3702 10280 3742 10600
rect 4062 10280 4102 10600
rect 3702 10240 4102 10280
rect 4714 10600 5114 10640
rect 4714 10280 4754 10600
rect 5074 10280 5114 10600
rect 4714 10240 5114 10280
rect 5726 10600 6126 10640
rect 5726 10280 5766 10600
rect 6086 10280 6126 10600
rect 5726 10240 6126 10280
rect 6738 10600 7138 10640
rect 6738 10280 6778 10600
rect 7098 10280 7138 10600
rect 6738 10240 7138 10280
rect -7430 9880 -7030 9920
rect -7430 9560 -7390 9880
rect -7070 9560 -7030 9880
rect -7430 9520 -7030 9560
rect -6418 9880 -6018 9920
rect -6418 9560 -6378 9880
rect -6058 9560 -6018 9880
rect -6418 9520 -6018 9560
rect -5406 9880 -5006 9920
rect -5406 9560 -5366 9880
rect -5046 9560 -5006 9880
rect -5406 9520 -5006 9560
rect -4394 9880 -3994 9920
rect -4394 9560 -4354 9880
rect -4034 9560 -3994 9880
rect -4394 9520 -3994 9560
rect -3382 9880 -2982 9920
rect -3382 9560 -3342 9880
rect -3022 9560 -2982 9880
rect -3382 9520 -2982 9560
rect -2370 9880 -1970 9920
rect -2370 9560 -2330 9880
rect -2010 9560 -1970 9880
rect -2370 9520 -1970 9560
rect -1358 9880 -958 9920
rect -1358 9560 -1318 9880
rect -998 9560 -958 9880
rect -1358 9520 -958 9560
rect -346 9880 54 9920
rect -346 9560 -306 9880
rect 14 9560 54 9880
rect -346 9520 54 9560
rect 666 9880 1066 9920
rect 666 9560 706 9880
rect 1026 9560 1066 9880
rect 666 9520 1066 9560
rect 1678 9880 2078 9920
rect 1678 9560 1718 9880
rect 2038 9560 2078 9880
rect 1678 9520 2078 9560
rect 2690 9880 3090 9920
rect 2690 9560 2730 9880
rect 3050 9560 3090 9880
rect 2690 9520 3090 9560
rect 3702 9880 4102 9920
rect 3702 9560 3742 9880
rect 4062 9560 4102 9880
rect 3702 9520 4102 9560
rect 4714 9880 5114 9920
rect 4714 9560 4754 9880
rect 5074 9560 5114 9880
rect 4714 9520 5114 9560
rect 5726 9880 6126 9920
rect 5726 9560 5766 9880
rect 6086 9560 6126 9880
rect 5726 9520 6126 9560
rect 6738 9880 7138 9920
rect 6738 9560 6778 9880
rect 7098 9560 7138 9880
rect 6738 9520 7138 9560
rect -7430 9160 -7030 9200
rect -7430 8840 -7390 9160
rect -7070 8840 -7030 9160
rect -7430 8800 -7030 8840
rect -6418 9160 -6018 9200
rect -6418 8840 -6378 9160
rect -6058 8840 -6018 9160
rect -6418 8800 -6018 8840
rect -5406 9160 -5006 9200
rect -5406 8840 -5366 9160
rect -5046 8840 -5006 9160
rect -5406 8800 -5006 8840
rect -4394 9160 -3994 9200
rect -4394 8840 -4354 9160
rect -4034 8840 -3994 9160
rect -4394 8800 -3994 8840
rect -3382 9160 -2982 9200
rect -3382 8840 -3342 9160
rect -3022 8840 -2982 9160
rect -3382 8800 -2982 8840
rect -2370 9160 -1970 9200
rect -2370 8840 -2330 9160
rect -2010 8840 -1970 9160
rect -2370 8800 -1970 8840
rect -1358 9160 -958 9200
rect -1358 8840 -1318 9160
rect -998 8840 -958 9160
rect -1358 8800 -958 8840
rect -346 9160 54 9200
rect -346 8840 -306 9160
rect 14 8840 54 9160
rect -346 8800 54 8840
rect 666 9160 1066 9200
rect 666 8840 706 9160
rect 1026 8840 1066 9160
rect 666 8800 1066 8840
rect 1678 9160 2078 9200
rect 1678 8840 1718 9160
rect 2038 8840 2078 9160
rect 1678 8800 2078 8840
rect 2690 9160 3090 9200
rect 2690 8840 2730 9160
rect 3050 8840 3090 9160
rect 2690 8800 3090 8840
rect 3702 9160 4102 9200
rect 3702 8840 3742 9160
rect 4062 8840 4102 9160
rect 3702 8800 4102 8840
rect 4714 9160 5114 9200
rect 4714 8840 4754 9160
rect 5074 8840 5114 9160
rect 4714 8800 5114 8840
rect 5726 9160 6126 9200
rect 5726 8840 5766 9160
rect 6086 8840 6126 9160
rect 5726 8800 6126 8840
rect 6738 9160 7138 9200
rect 6738 8840 6778 9160
rect 7098 8840 7138 9160
rect 6738 8800 7138 8840
rect -7430 8440 -7030 8480
rect -7430 8120 -7390 8440
rect -7070 8120 -7030 8440
rect -7430 8080 -7030 8120
rect -6418 8440 -6018 8480
rect -6418 8120 -6378 8440
rect -6058 8120 -6018 8440
rect -6418 8080 -6018 8120
rect -5406 8440 -5006 8480
rect -5406 8120 -5366 8440
rect -5046 8120 -5006 8440
rect -5406 8080 -5006 8120
rect -4394 8440 -3994 8480
rect -4394 8120 -4354 8440
rect -4034 8120 -3994 8440
rect -4394 8080 -3994 8120
rect -3382 8440 -2982 8480
rect -3382 8120 -3342 8440
rect -3022 8120 -2982 8440
rect -3382 8080 -2982 8120
rect -2370 8440 -1970 8480
rect -2370 8120 -2330 8440
rect -2010 8120 -1970 8440
rect -2370 8080 -1970 8120
rect -1358 8440 -958 8480
rect -1358 8120 -1318 8440
rect -998 8120 -958 8440
rect -1358 8080 -958 8120
rect -346 8440 54 8480
rect -346 8120 -306 8440
rect 14 8120 54 8440
rect -346 8080 54 8120
rect 666 8440 1066 8480
rect 666 8120 706 8440
rect 1026 8120 1066 8440
rect 666 8080 1066 8120
rect 1678 8440 2078 8480
rect 1678 8120 1718 8440
rect 2038 8120 2078 8440
rect 1678 8080 2078 8120
rect 2690 8440 3090 8480
rect 2690 8120 2730 8440
rect 3050 8120 3090 8440
rect 2690 8080 3090 8120
rect 3702 8440 4102 8480
rect 3702 8120 3742 8440
rect 4062 8120 4102 8440
rect 3702 8080 4102 8120
rect 4714 8440 5114 8480
rect 4714 8120 4754 8440
rect 5074 8120 5114 8440
rect 4714 8080 5114 8120
rect 5726 8440 6126 8480
rect 5726 8120 5766 8440
rect 6086 8120 6126 8440
rect 5726 8080 6126 8120
rect 6738 8440 7138 8480
rect 6738 8120 6778 8440
rect 7098 8120 7138 8440
rect 6738 8080 7138 8120
rect -7430 7720 -7030 7760
rect -7430 7400 -7390 7720
rect -7070 7400 -7030 7720
rect -7430 7360 -7030 7400
rect -6418 7720 -6018 7760
rect -6418 7400 -6378 7720
rect -6058 7400 -6018 7720
rect -6418 7360 -6018 7400
rect -5406 7720 -5006 7760
rect -5406 7400 -5366 7720
rect -5046 7400 -5006 7720
rect -5406 7360 -5006 7400
rect -4394 7720 -3994 7760
rect -4394 7400 -4354 7720
rect -4034 7400 -3994 7720
rect -4394 7360 -3994 7400
rect -3382 7720 -2982 7760
rect -3382 7400 -3342 7720
rect -3022 7400 -2982 7720
rect -3382 7360 -2982 7400
rect -2370 7720 -1970 7760
rect -2370 7400 -2330 7720
rect -2010 7400 -1970 7720
rect -2370 7360 -1970 7400
rect -1358 7720 -958 7760
rect -1358 7400 -1318 7720
rect -998 7400 -958 7720
rect -1358 7360 -958 7400
rect -346 7720 54 7760
rect -346 7400 -306 7720
rect 14 7400 54 7720
rect -346 7360 54 7400
rect 666 7720 1066 7760
rect 666 7400 706 7720
rect 1026 7400 1066 7720
rect 666 7360 1066 7400
rect 1678 7720 2078 7760
rect 1678 7400 1718 7720
rect 2038 7400 2078 7720
rect 1678 7360 2078 7400
rect 2690 7720 3090 7760
rect 2690 7400 2730 7720
rect 3050 7400 3090 7720
rect 2690 7360 3090 7400
rect 3702 7720 4102 7760
rect 3702 7400 3742 7720
rect 4062 7400 4102 7720
rect 3702 7360 4102 7400
rect 4714 7720 5114 7760
rect 4714 7400 4754 7720
rect 5074 7400 5114 7720
rect 4714 7360 5114 7400
rect 5726 7720 6126 7760
rect 5726 7400 5766 7720
rect 6086 7400 6126 7720
rect 5726 7360 6126 7400
rect 6738 7720 7138 7760
rect 6738 7400 6778 7720
rect 7098 7400 7138 7720
rect 6738 7360 7138 7400
rect -7430 7000 -7030 7040
rect -7430 6680 -7390 7000
rect -7070 6680 -7030 7000
rect -7430 6640 -7030 6680
rect -6418 7000 -6018 7040
rect -6418 6680 -6378 7000
rect -6058 6680 -6018 7000
rect -6418 6640 -6018 6680
rect -5406 7000 -5006 7040
rect -5406 6680 -5366 7000
rect -5046 6680 -5006 7000
rect -5406 6640 -5006 6680
rect -4394 7000 -3994 7040
rect -4394 6680 -4354 7000
rect -4034 6680 -3994 7000
rect -4394 6640 -3994 6680
rect -3382 7000 -2982 7040
rect -3382 6680 -3342 7000
rect -3022 6680 -2982 7000
rect -3382 6640 -2982 6680
rect -2370 7000 -1970 7040
rect -2370 6680 -2330 7000
rect -2010 6680 -1970 7000
rect -2370 6640 -1970 6680
rect -1358 7000 -958 7040
rect -1358 6680 -1318 7000
rect -998 6680 -958 7000
rect -1358 6640 -958 6680
rect -346 7000 54 7040
rect -346 6680 -306 7000
rect 14 6680 54 7000
rect -346 6640 54 6680
rect 666 7000 1066 7040
rect 666 6680 706 7000
rect 1026 6680 1066 7000
rect 666 6640 1066 6680
rect 1678 7000 2078 7040
rect 1678 6680 1718 7000
rect 2038 6680 2078 7000
rect 1678 6640 2078 6680
rect 2690 7000 3090 7040
rect 2690 6680 2730 7000
rect 3050 6680 3090 7000
rect 2690 6640 3090 6680
rect 3702 7000 4102 7040
rect 3702 6680 3742 7000
rect 4062 6680 4102 7000
rect 3702 6640 4102 6680
rect 4714 7000 5114 7040
rect 4714 6680 4754 7000
rect 5074 6680 5114 7000
rect 4714 6640 5114 6680
rect 5726 7000 6126 7040
rect 5726 6680 5766 7000
rect 6086 6680 6126 7000
rect 5726 6640 6126 6680
rect 6738 7000 7138 7040
rect 6738 6680 6778 7000
rect 7098 6680 7138 7000
rect 6738 6640 7138 6680
rect -7430 6280 -7030 6320
rect -7430 5960 -7390 6280
rect -7070 5960 -7030 6280
rect -7430 5920 -7030 5960
rect -6418 6280 -6018 6320
rect -6418 5960 -6378 6280
rect -6058 5960 -6018 6280
rect -6418 5920 -6018 5960
rect -5406 6280 -5006 6320
rect -5406 5960 -5366 6280
rect -5046 5960 -5006 6280
rect -5406 5920 -5006 5960
rect -4394 6280 -3994 6320
rect -4394 5960 -4354 6280
rect -4034 5960 -3994 6280
rect -4394 5920 -3994 5960
rect -3382 6280 -2982 6320
rect -3382 5960 -3342 6280
rect -3022 5960 -2982 6280
rect -3382 5920 -2982 5960
rect -2370 6280 -1970 6320
rect -2370 5960 -2330 6280
rect -2010 5960 -1970 6280
rect -2370 5920 -1970 5960
rect -1358 6280 -958 6320
rect -1358 5960 -1318 6280
rect -998 5960 -958 6280
rect -1358 5920 -958 5960
rect -346 6280 54 6320
rect -346 5960 -306 6280
rect 14 5960 54 6280
rect -346 5920 54 5960
rect 666 6280 1066 6320
rect 666 5960 706 6280
rect 1026 5960 1066 6280
rect 666 5920 1066 5960
rect 1678 6280 2078 6320
rect 1678 5960 1718 6280
rect 2038 5960 2078 6280
rect 1678 5920 2078 5960
rect 2690 6280 3090 6320
rect 2690 5960 2730 6280
rect 3050 5960 3090 6280
rect 2690 5920 3090 5960
rect 3702 6280 4102 6320
rect 3702 5960 3742 6280
rect 4062 5960 4102 6280
rect 3702 5920 4102 5960
rect 4714 6280 5114 6320
rect 4714 5960 4754 6280
rect 5074 5960 5114 6280
rect 4714 5920 5114 5960
rect 5726 6280 6126 6320
rect 5726 5960 5766 6280
rect 6086 5960 6126 6280
rect 5726 5920 6126 5960
rect 6738 6280 7138 6320
rect 6738 5960 6778 6280
rect 7098 5960 7138 6280
rect 6738 5920 7138 5960
rect -7430 5560 -7030 5600
rect -7430 5240 -7390 5560
rect -7070 5240 -7030 5560
rect -7430 5200 -7030 5240
rect -6418 5560 -6018 5600
rect -6418 5240 -6378 5560
rect -6058 5240 -6018 5560
rect -6418 5200 -6018 5240
rect -5406 5560 -5006 5600
rect -5406 5240 -5366 5560
rect -5046 5240 -5006 5560
rect -5406 5200 -5006 5240
rect -4394 5560 -3994 5600
rect -4394 5240 -4354 5560
rect -4034 5240 -3994 5560
rect -4394 5200 -3994 5240
rect -3382 5560 -2982 5600
rect -3382 5240 -3342 5560
rect -3022 5240 -2982 5560
rect -3382 5200 -2982 5240
rect -2370 5560 -1970 5600
rect -2370 5240 -2330 5560
rect -2010 5240 -1970 5560
rect -2370 5200 -1970 5240
rect -1358 5560 -958 5600
rect -1358 5240 -1318 5560
rect -998 5240 -958 5560
rect -1358 5200 -958 5240
rect -346 5560 54 5600
rect -346 5240 -306 5560
rect 14 5240 54 5560
rect -346 5200 54 5240
rect 666 5560 1066 5600
rect 666 5240 706 5560
rect 1026 5240 1066 5560
rect 666 5200 1066 5240
rect 1678 5560 2078 5600
rect 1678 5240 1718 5560
rect 2038 5240 2078 5560
rect 1678 5200 2078 5240
rect 2690 5560 3090 5600
rect 2690 5240 2730 5560
rect 3050 5240 3090 5560
rect 2690 5200 3090 5240
rect 3702 5560 4102 5600
rect 3702 5240 3742 5560
rect 4062 5240 4102 5560
rect 3702 5200 4102 5240
rect 4714 5560 5114 5600
rect 4714 5240 4754 5560
rect 5074 5240 5114 5560
rect 4714 5200 5114 5240
rect 5726 5560 6126 5600
rect 5726 5240 5766 5560
rect 6086 5240 6126 5560
rect 5726 5200 6126 5240
rect 6738 5560 7138 5600
rect 6738 5240 6778 5560
rect 7098 5240 7138 5560
rect 6738 5200 7138 5240
rect -7430 4840 -7030 4880
rect -7430 4520 -7390 4840
rect -7070 4520 -7030 4840
rect -7430 4480 -7030 4520
rect -6418 4840 -6018 4880
rect -6418 4520 -6378 4840
rect -6058 4520 -6018 4840
rect -6418 4480 -6018 4520
rect -5406 4840 -5006 4880
rect -5406 4520 -5366 4840
rect -5046 4520 -5006 4840
rect -5406 4480 -5006 4520
rect -4394 4840 -3994 4880
rect -4394 4520 -4354 4840
rect -4034 4520 -3994 4840
rect -4394 4480 -3994 4520
rect -3382 4840 -2982 4880
rect -3382 4520 -3342 4840
rect -3022 4520 -2982 4840
rect -3382 4480 -2982 4520
rect -2370 4840 -1970 4880
rect -2370 4520 -2330 4840
rect -2010 4520 -1970 4840
rect -2370 4480 -1970 4520
rect -1358 4840 -958 4880
rect -1358 4520 -1318 4840
rect -998 4520 -958 4840
rect -1358 4480 -958 4520
rect -346 4840 54 4880
rect -346 4520 -306 4840
rect 14 4520 54 4840
rect -346 4480 54 4520
rect 666 4840 1066 4880
rect 666 4520 706 4840
rect 1026 4520 1066 4840
rect 666 4480 1066 4520
rect 1678 4840 2078 4880
rect 1678 4520 1718 4840
rect 2038 4520 2078 4840
rect 1678 4480 2078 4520
rect 2690 4840 3090 4880
rect 2690 4520 2730 4840
rect 3050 4520 3090 4840
rect 2690 4480 3090 4520
rect 3702 4840 4102 4880
rect 3702 4520 3742 4840
rect 4062 4520 4102 4840
rect 3702 4480 4102 4520
rect 4714 4840 5114 4880
rect 4714 4520 4754 4840
rect 5074 4520 5114 4840
rect 4714 4480 5114 4520
rect 5726 4840 6126 4880
rect 5726 4520 5766 4840
rect 6086 4520 6126 4840
rect 5726 4480 6126 4520
rect 6738 4840 7138 4880
rect 6738 4520 6778 4840
rect 7098 4520 7138 4840
rect 6738 4480 7138 4520
rect -7430 4120 -7030 4160
rect -7430 3800 -7390 4120
rect -7070 3800 -7030 4120
rect -7430 3760 -7030 3800
rect -6418 4120 -6018 4160
rect -6418 3800 -6378 4120
rect -6058 3800 -6018 4120
rect -6418 3760 -6018 3800
rect -5406 4120 -5006 4160
rect -5406 3800 -5366 4120
rect -5046 3800 -5006 4120
rect -5406 3760 -5006 3800
rect -4394 4120 -3994 4160
rect -4394 3800 -4354 4120
rect -4034 3800 -3994 4120
rect -4394 3760 -3994 3800
rect -3382 4120 -2982 4160
rect -3382 3800 -3342 4120
rect -3022 3800 -2982 4120
rect -3382 3760 -2982 3800
rect -2370 4120 -1970 4160
rect -2370 3800 -2330 4120
rect -2010 3800 -1970 4120
rect -2370 3760 -1970 3800
rect -1358 4120 -958 4160
rect -1358 3800 -1318 4120
rect -998 3800 -958 4120
rect -1358 3760 -958 3800
rect -346 4120 54 4160
rect -346 3800 -306 4120
rect 14 3800 54 4120
rect -346 3760 54 3800
rect 666 4120 1066 4160
rect 666 3800 706 4120
rect 1026 3800 1066 4120
rect 666 3760 1066 3800
rect 1678 4120 2078 4160
rect 1678 3800 1718 4120
rect 2038 3800 2078 4120
rect 1678 3760 2078 3800
rect 2690 4120 3090 4160
rect 2690 3800 2730 4120
rect 3050 3800 3090 4120
rect 2690 3760 3090 3800
rect 3702 4120 4102 4160
rect 3702 3800 3742 4120
rect 4062 3800 4102 4120
rect 3702 3760 4102 3800
rect 4714 4120 5114 4160
rect 4714 3800 4754 4120
rect 5074 3800 5114 4120
rect 4714 3760 5114 3800
rect 5726 4120 6126 4160
rect 5726 3800 5766 4120
rect 6086 3800 6126 4120
rect 5726 3760 6126 3800
rect 6738 4120 7138 4160
rect 6738 3800 6778 4120
rect 7098 3800 7138 4120
rect 6738 3760 7138 3800
rect -7430 3400 -7030 3440
rect -7430 3080 -7390 3400
rect -7070 3080 -7030 3400
rect -7430 3040 -7030 3080
rect -6418 3400 -6018 3440
rect -6418 3080 -6378 3400
rect -6058 3080 -6018 3400
rect -6418 3040 -6018 3080
rect -5406 3400 -5006 3440
rect -5406 3080 -5366 3400
rect -5046 3080 -5006 3400
rect -5406 3040 -5006 3080
rect -4394 3400 -3994 3440
rect -4394 3080 -4354 3400
rect -4034 3080 -3994 3400
rect -4394 3040 -3994 3080
rect -3382 3400 -2982 3440
rect -3382 3080 -3342 3400
rect -3022 3080 -2982 3400
rect -3382 3040 -2982 3080
rect -2370 3400 -1970 3440
rect -2370 3080 -2330 3400
rect -2010 3080 -1970 3400
rect -2370 3040 -1970 3080
rect -1358 3400 -958 3440
rect -1358 3080 -1318 3400
rect -998 3080 -958 3400
rect -1358 3040 -958 3080
rect -346 3400 54 3440
rect -346 3080 -306 3400
rect 14 3080 54 3400
rect -346 3040 54 3080
rect 666 3400 1066 3440
rect 666 3080 706 3400
rect 1026 3080 1066 3400
rect 666 3040 1066 3080
rect 1678 3400 2078 3440
rect 1678 3080 1718 3400
rect 2038 3080 2078 3400
rect 1678 3040 2078 3080
rect 2690 3400 3090 3440
rect 2690 3080 2730 3400
rect 3050 3080 3090 3400
rect 2690 3040 3090 3080
rect 3702 3400 4102 3440
rect 3702 3080 3742 3400
rect 4062 3080 4102 3400
rect 3702 3040 4102 3080
rect 4714 3400 5114 3440
rect 4714 3080 4754 3400
rect 5074 3080 5114 3400
rect 4714 3040 5114 3080
rect 5726 3400 6126 3440
rect 5726 3080 5766 3400
rect 6086 3080 6126 3400
rect 5726 3040 6126 3080
rect 6738 3400 7138 3440
rect 6738 3080 6778 3400
rect 7098 3080 7138 3400
rect 6738 3040 7138 3080
rect -7430 2680 -7030 2720
rect -7430 2360 -7390 2680
rect -7070 2360 -7030 2680
rect -7430 2320 -7030 2360
rect -6418 2680 -6018 2720
rect -6418 2360 -6378 2680
rect -6058 2360 -6018 2680
rect -6418 2320 -6018 2360
rect -5406 2680 -5006 2720
rect -5406 2360 -5366 2680
rect -5046 2360 -5006 2680
rect -5406 2320 -5006 2360
rect -4394 2680 -3994 2720
rect -4394 2360 -4354 2680
rect -4034 2360 -3994 2680
rect -4394 2320 -3994 2360
rect -3382 2680 -2982 2720
rect -3382 2360 -3342 2680
rect -3022 2360 -2982 2680
rect -3382 2320 -2982 2360
rect -2370 2680 -1970 2720
rect -2370 2360 -2330 2680
rect -2010 2360 -1970 2680
rect -2370 2320 -1970 2360
rect -1358 2680 -958 2720
rect -1358 2360 -1318 2680
rect -998 2360 -958 2680
rect -1358 2320 -958 2360
rect -346 2680 54 2720
rect -346 2360 -306 2680
rect 14 2360 54 2680
rect -346 2320 54 2360
rect 666 2680 1066 2720
rect 666 2360 706 2680
rect 1026 2360 1066 2680
rect 666 2320 1066 2360
rect 1678 2680 2078 2720
rect 1678 2360 1718 2680
rect 2038 2360 2078 2680
rect 1678 2320 2078 2360
rect 2690 2680 3090 2720
rect 2690 2360 2730 2680
rect 3050 2360 3090 2680
rect 2690 2320 3090 2360
rect 3702 2680 4102 2720
rect 3702 2360 3742 2680
rect 4062 2360 4102 2680
rect 3702 2320 4102 2360
rect 4714 2680 5114 2720
rect 4714 2360 4754 2680
rect 5074 2360 5114 2680
rect 4714 2320 5114 2360
rect 5726 2680 6126 2720
rect 5726 2360 5766 2680
rect 6086 2360 6126 2680
rect 5726 2320 6126 2360
rect 6738 2680 7138 2720
rect 6738 2360 6778 2680
rect 7098 2360 7138 2680
rect 6738 2320 7138 2360
rect -7430 1960 -7030 2000
rect -7430 1640 -7390 1960
rect -7070 1640 -7030 1960
rect -7430 1600 -7030 1640
rect -6418 1960 -6018 2000
rect -6418 1640 -6378 1960
rect -6058 1640 -6018 1960
rect -6418 1600 -6018 1640
rect -5406 1960 -5006 2000
rect -5406 1640 -5366 1960
rect -5046 1640 -5006 1960
rect -5406 1600 -5006 1640
rect -4394 1960 -3994 2000
rect -4394 1640 -4354 1960
rect -4034 1640 -3994 1960
rect -4394 1600 -3994 1640
rect -3382 1960 -2982 2000
rect -3382 1640 -3342 1960
rect -3022 1640 -2982 1960
rect -3382 1600 -2982 1640
rect -2370 1960 -1970 2000
rect -2370 1640 -2330 1960
rect -2010 1640 -1970 1960
rect -2370 1600 -1970 1640
rect -1358 1960 -958 2000
rect -1358 1640 -1318 1960
rect -998 1640 -958 1960
rect -1358 1600 -958 1640
rect -346 1960 54 2000
rect -346 1640 -306 1960
rect 14 1640 54 1960
rect -346 1600 54 1640
rect 666 1960 1066 2000
rect 666 1640 706 1960
rect 1026 1640 1066 1960
rect 666 1600 1066 1640
rect 1678 1960 2078 2000
rect 1678 1640 1718 1960
rect 2038 1640 2078 1960
rect 1678 1600 2078 1640
rect 2690 1960 3090 2000
rect 2690 1640 2730 1960
rect 3050 1640 3090 1960
rect 2690 1600 3090 1640
rect 3702 1960 4102 2000
rect 3702 1640 3742 1960
rect 4062 1640 4102 1960
rect 3702 1600 4102 1640
rect 4714 1960 5114 2000
rect 4714 1640 4754 1960
rect 5074 1640 5114 1960
rect 4714 1600 5114 1640
rect 5726 1960 6126 2000
rect 5726 1640 5766 1960
rect 6086 1640 6126 1960
rect 5726 1600 6126 1640
rect 6738 1960 7138 2000
rect 6738 1640 6778 1960
rect 7098 1640 7138 1960
rect 6738 1600 7138 1640
rect -7430 1240 -7030 1280
rect -7430 920 -7390 1240
rect -7070 920 -7030 1240
rect -7430 880 -7030 920
rect -6418 1240 -6018 1280
rect -6418 920 -6378 1240
rect -6058 920 -6018 1240
rect -6418 880 -6018 920
rect -5406 1240 -5006 1280
rect -5406 920 -5366 1240
rect -5046 920 -5006 1240
rect -5406 880 -5006 920
rect -4394 1240 -3994 1280
rect -4394 920 -4354 1240
rect -4034 920 -3994 1240
rect -4394 880 -3994 920
rect -3382 1240 -2982 1280
rect -3382 920 -3342 1240
rect -3022 920 -2982 1240
rect -3382 880 -2982 920
rect -2370 1240 -1970 1280
rect -2370 920 -2330 1240
rect -2010 920 -1970 1240
rect -2370 880 -1970 920
rect -1358 1240 -958 1280
rect -1358 920 -1318 1240
rect -998 920 -958 1240
rect -1358 880 -958 920
rect -346 1240 54 1280
rect -346 920 -306 1240
rect 14 920 54 1240
rect -346 880 54 920
rect 666 1240 1066 1280
rect 666 920 706 1240
rect 1026 920 1066 1240
rect 666 880 1066 920
rect 1678 1240 2078 1280
rect 1678 920 1718 1240
rect 2038 920 2078 1240
rect 1678 880 2078 920
rect 2690 1240 3090 1280
rect 2690 920 2730 1240
rect 3050 920 3090 1240
rect 2690 880 3090 920
rect 3702 1240 4102 1280
rect 3702 920 3742 1240
rect 4062 920 4102 1240
rect 3702 880 4102 920
rect 4714 1240 5114 1280
rect 4714 920 4754 1240
rect 5074 920 5114 1240
rect 4714 880 5114 920
rect 5726 1240 6126 1280
rect 5726 920 5766 1240
rect 6086 920 6126 1240
rect 5726 880 6126 920
rect 6738 1240 7138 1280
rect 6738 920 6778 1240
rect 7098 920 7138 1240
rect 6738 880 7138 920
rect -7430 520 -7030 560
rect -7430 200 -7390 520
rect -7070 200 -7030 520
rect -7430 160 -7030 200
rect -6418 520 -6018 560
rect -6418 200 -6378 520
rect -6058 200 -6018 520
rect -6418 160 -6018 200
rect -5406 520 -5006 560
rect -5406 200 -5366 520
rect -5046 200 -5006 520
rect -5406 160 -5006 200
rect -4394 520 -3994 560
rect -4394 200 -4354 520
rect -4034 200 -3994 520
rect -4394 160 -3994 200
rect -3382 520 -2982 560
rect -3382 200 -3342 520
rect -3022 200 -2982 520
rect -3382 160 -2982 200
rect -2370 520 -1970 560
rect -2370 200 -2330 520
rect -2010 200 -1970 520
rect -2370 160 -1970 200
rect -1358 520 -958 560
rect -1358 200 -1318 520
rect -998 200 -958 520
rect -1358 160 -958 200
rect -346 520 54 560
rect -346 200 -306 520
rect 14 200 54 520
rect -346 160 54 200
rect 666 520 1066 560
rect 666 200 706 520
rect 1026 200 1066 520
rect 666 160 1066 200
rect 1678 520 2078 560
rect 1678 200 1718 520
rect 2038 200 2078 520
rect 1678 160 2078 200
rect 2690 520 3090 560
rect 2690 200 2730 520
rect 3050 200 3090 520
rect 2690 160 3090 200
rect 3702 520 4102 560
rect 3702 200 3742 520
rect 4062 200 4102 520
rect 3702 160 4102 200
rect 4714 520 5114 560
rect 4714 200 4754 520
rect 5074 200 5114 520
rect 4714 160 5114 200
rect 5726 520 6126 560
rect 5726 200 5766 520
rect 6086 200 6126 520
rect 5726 160 6126 200
rect 6738 520 7138 560
rect 6738 200 6778 520
rect 7098 200 7138 520
rect 6738 160 7138 200
rect -7430 -200 -7030 -160
rect -7430 -520 -7390 -200
rect -7070 -520 -7030 -200
rect -7430 -560 -7030 -520
rect -6418 -200 -6018 -160
rect -6418 -520 -6378 -200
rect -6058 -520 -6018 -200
rect -6418 -560 -6018 -520
rect -5406 -200 -5006 -160
rect -5406 -520 -5366 -200
rect -5046 -520 -5006 -200
rect -5406 -560 -5006 -520
rect -4394 -200 -3994 -160
rect -4394 -520 -4354 -200
rect -4034 -520 -3994 -200
rect -4394 -560 -3994 -520
rect -3382 -200 -2982 -160
rect -3382 -520 -3342 -200
rect -3022 -520 -2982 -200
rect -3382 -560 -2982 -520
rect -2370 -200 -1970 -160
rect -2370 -520 -2330 -200
rect -2010 -520 -1970 -200
rect -2370 -560 -1970 -520
rect -1358 -200 -958 -160
rect -1358 -520 -1318 -200
rect -998 -520 -958 -200
rect -1358 -560 -958 -520
rect -346 -200 54 -160
rect -346 -520 -306 -200
rect 14 -520 54 -200
rect -346 -560 54 -520
rect 666 -200 1066 -160
rect 666 -520 706 -200
rect 1026 -520 1066 -200
rect 666 -560 1066 -520
rect 1678 -200 2078 -160
rect 1678 -520 1718 -200
rect 2038 -520 2078 -200
rect 1678 -560 2078 -520
rect 2690 -200 3090 -160
rect 2690 -520 2730 -200
rect 3050 -520 3090 -200
rect 2690 -560 3090 -520
rect 3702 -200 4102 -160
rect 3702 -520 3742 -200
rect 4062 -520 4102 -200
rect 3702 -560 4102 -520
rect 4714 -200 5114 -160
rect 4714 -520 4754 -200
rect 5074 -520 5114 -200
rect 4714 -560 5114 -520
rect 5726 -200 6126 -160
rect 5726 -520 5766 -200
rect 6086 -520 6126 -200
rect 5726 -560 6126 -520
rect 6738 -200 7138 -160
rect 6738 -520 6778 -200
rect 7098 -520 7138 -200
rect 6738 -560 7138 -520
rect -7430 -920 -7030 -880
rect -7430 -1240 -7390 -920
rect -7070 -1240 -7030 -920
rect -7430 -1280 -7030 -1240
rect -6418 -920 -6018 -880
rect -6418 -1240 -6378 -920
rect -6058 -1240 -6018 -920
rect -6418 -1280 -6018 -1240
rect -5406 -920 -5006 -880
rect -5406 -1240 -5366 -920
rect -5046 -1240 -5006 -920
rect -5406 -1280 -5006 -1240
rect -4394 -920 -3994 -880
rect -4394 -1240 -4354 -920
rect -4034 -1240 -3994 -920
rect -4394 -1280 -3994 -1240
rect -3382 -920 -2982 -880
rect -3382 -1240 -3342 -920
rect -3022 -1240 -2982 -920
rect -3382 -1280 -2982 -1240
rect -2370 -920 -1970 -880
rect -2370 -1240 -2330 -920
rect -2010 -1240 -1970 -920
rect -2370 -1280 -1970 -1240
rect -1358 -920 -958 -880
rect -1358 -1240 -1318 -920
rect -998 -1240 -958 -920
rect -1358 -1280 -958 -1240
rect -346 -920 54 -880
rect -346 -1240 -306 -920
rect 14 -1240 54 -920
rect -346 -1280 54 -1240
rect 666 -920 1066 -880
rect 666 -1240 706 -920
rect 1026 -1240 1066 -920
rect 666 -1280 1066 -1240
rect 1678 -920 2078 -880
rect 1678 -1240 1718 -920
rect 2038 -1240 2078 -920
rect 1678 -1280 2078 -1240
rect 2690 -920 3090 -880
rect 2690 -1240 2730 -920
rect 3050 -1240 3090 -920
rect 2690 -1280 3090 -1240
rect 3702 -920 4102 -880
rect 3702 -1240 3742 -920
rect 4062 -1240 4102 -920
rect 3702 -1280 4102 -1240
rect 4714 -920 5114 -880
rect 4714 -1240 4754 -920
rect 5074 -1240 5114 -920
rect 4714 -1280 5114 -1240
rect 5726 -920 6126 -880
rect 5726 -1240 5766 -920
rect 6086 -1240 6126 -920
rect 5726 -1280 6126 -1240
rect 6738 -920 7138 -880
rect 6738 -1240 6778 -920
rect 7098 -1240 7138 -920
rect 6738 -1280 7138 -1240
rect -7430 -1640 -7030 -1600
rect -7430 -1960 -7390 -1640
rect -7070 -1960 -7030 -1640
rect -7430 -2000 -7030 -1960
rect -6418 -1640 -6018 -1600
rect -6418 -1960 -6378 -1640
rect -6058 -1960 -6018 -1640
rect -6418 -2000 -6018 -1960
rect -5406 -1640 -5006 -1600
rect -5406 -1960 -5366 -1640
rect -5046 -1960 -5006 -1640
rect -5406 -2000 -5006 -1960
rect -4394 -1640 -3994 -1600
rect -4394 -1960 -4354 -1640
rect -4034 -1960 -3994 -1640
rect -4394 -2000 -3994 -1960
rect -3382 -1640 -2982 -1600
rect -3382 -1960 -3342 -1640
rect -3022 -1960 -2982 -1640
rect -3382 -2000 -2982 -1960
rect -2370 -1640 -1970 -1600
rect -2370 -1960 -2330 -1640
rect -2010 -1960 -1970 -1640
rect -2370 -2000 -1970 -1960
rect -1358 -1640 -958 -1600
rect -1358 -1960 -1318 -1640
rect -998 -1960 -958 -1640
rect -1358 -2000 -958 -1960
rect -346 -1640 54 -1600
rect -346 -1960 -306 -1640
rect 14 -1960 54 -1640
rect -346 -2000 54 -1960
rect 666 -1640 1066 -1600
rect 666 -1960 706 -1640
rect 1026 -1960 1066 -1640
rect 666 -2000 1066 -1960
rect 1678 -1640 2078 -1600
rect 1678 -1960 1718 -1640
rect 2038 -1960 2078 -1640
rect 1678 -2000 2078 -1960
rect 2690 -1640 3090 -1600
rect 2690 -1960 2730 -1640
rect 3050 -1960 3090 -1640
rect 2690 -2000 3090 -1960
rect 3702 -1640 4102 -1600
rect 3702 -1960 3742 -1640
rect 4062 -1960 4102 -1640
rect 3702 -2000 4102 -1960
rect 4714 -1640 5114 -1600
rect 4714 -1960 4754 -1640
rect 5074 -1960 5114 -1640
rect 4714 -2000 5114 -1960
rect 5726 -1640 6126 -1600
rect 5726 -1960 5766 -1640
rect 6086 -1960 6126 -1640
rect 5726 -2000 6126 -1960
rect 6738 -1640 7138 -1600
rect 6738 -1960 6778 -1640
rect 7098 -1960 7138 -1640
rect 6738 -2000 7138 -1960
rect -7430 -2360 -7030 -2320
rect -7430 -2680 -7390 -2360
rect -7070 -2680 -7030 -2360
rect -7430 -2720 -7030 -2680
rect -6418 -2360 -6018 -2320
rect -6418 -2680 -6378 -2360
rect -6058 -2680 -6018 -2360
rect -6418 -2720 -6018 -2680
rect -5406 -2360 -5006 -2320
rect -5406 -2680 -5366 -2360
rect -5046 -2680 -5006 -2360
rect -5406 -2720 -5006 -2680
rect -4394 -2360 -3994 -2320
rect -4394 -2680 -4354 -2360
rect -4034 -2680 -3994 -2360
rect -4394 -2720 -3994 -2680
rect -3382 -2360 -2982 -2320
rect -3382 -2680 -3342 -2360
rect -3022 -2680 -2982 -2360
rect -3382 -2720 -2982 -2680
rect -2370 -2360 -1970 -2320
rect -2370 -2680 -2330 -2360
rect -2010 -2680 -1970 -2360
rect -2370 -2720 -1970 -2680
rect -1358 -2360 -958 -2320
rect -1358 -2680 -1318 -2360
rect -998 -2680 -958 -2360
rect -1358 -2720 -958 -2680
rect -346 -2360 54 -2320
rect -346 -2680 -306 -2360
rect 14 -2680 54 -2360
rect -346 -2720 54 -2680
rect 666 -2360 1066 -2320
rect 666 -2680 706 -2360
rect 1026 -2680 1066 -2360
rect 666 -2720 1066 -2680
rect 1678 -2360 2078 -2320
rect 1678 -2680 1718 -2360
rect 2038 -2680 2078 -2360
rect 1678 -2720 2078 -2680
rect 2690 -2360 3090 -2320
rect 2690 -2680 2730 -2360
rect 3050 -2680 3090 -2360
rect 2690 -2720 3090 -2680
rect 3702 -2360 4102 -2320
rect 3702 -2680 3742 -2360
rect 4062 -2680 4102 -2360
rect 3702 -2720 4102 -2680
rect 4714 -2360 5114 -2320
rect 4714 -2680 4754 -2360
rect 5074 -2680 5114 -2360
rect 4714 -2720 5114 -2680
rect 5726 -2360 6126 -2320
rect 5726 -2680 5766 -2360
rect 6086 -2680 6126 -2360
rect 5726 -2720 6126 -2680
rect 6738 -2360 7138 -2320
rect 6738 -2680 6778 -2360
rect 7098 -2680 7138 -2360
rect 6738 -2720 7138 -2680
rect -7430 -3080 -7030 -3040
rect -7430 -3400 -7390 -3080
rect -7070 -3400 -7030 -3080
rect -7430 -3440 -7030 -3400
rect -6418 -3080 -6018 -3040
rect -6418 -3400 -6378 -3080
rect -6058 -3400 -6018 -3080
rect -6418 -3440 -6018 -3400
rect -5406 -3080 -5006 -3040
rect -5406 -3400 -5366 -3080
rect -5046 -3400 -5006 -3080
rect -5406 -3440 -5006 -3400
rect -4394 -3080 -3994 -3040
rect -4394 -3400 -4354 -3080
rect -4034 -3400 -3994 -3080
rect -4394 -3440 -3994 -3400
rect -3382 -3080 -2982 -3040
rect -3382 -3400 -3342 -3080
rect -3022 -3400 -2982 -3080
rect -3382 -3440 -2982 -3400
rect -2370 -3080 -1970 -3040
rect -2370 -3400 -2330 -3080
rect -2010 -3400 -1970 -3080
rect -2370 -3440 -1970 -3400
rect -1358 -3080 -958 -3040
rect -1358 -3400 -1318 -3080
rect -998 -3400 -958 -3080
rect -1358 -3440 -958 -3400
rect -346 -3080 54 -3040
rect -346 -3400 -306 -3080
rect 14 -3400 54 -3080
rect -346 -3440 54 -3400
rect 666 -3080 1066 -3040
rect 666 -3400 706 -3080
rect 1026 -3400 1066 -3080
rect 666 -3440 1066 -3400
rect 1678 -3080 2078 -3040
rect 1678 -3400 1718 -3080
rect 2038 -3400 2078 -3080
rect 1678 -3440 2078 -3400
rect 2690 -3080 3090 -3040
rect 2690 -3400 2730 -3080
rect 3050 -3400 3090 -3080
rect 2690 -3440 3090 -3400
rect 3702 -3080 4102 -3040
rect 3702 -3400 3742 -3080
rect 4062 -3400 4102 -3080
rect 3702 -3440 4102 -3400
rect 4714 -3080 5114 -3040
rect 4714 -3400 4754 -3080
rect 5074 -3400 5114 -3080
rect 4714 -3440 5114 -3400
rect 5726 -3080 6126 -3040
rect 5726 -3400 5766 -3080
rect 6086 -3400 6126 -3080
rect 5726 -3440 6126 -3400
rect 6738 -3080 7138 -3040
rect 6738 -3400 6778 -3080
rect 7098 -3400 7138 -3080
rect 6738 -3440 7138 -3400
rect -7430 -3800 -7030 -3760
rect -7430 -4120 -7390 -3800
rect -7070 -4120 -7030 -3800
rect -7430 -4160 -7030 -4120
rect -6418 -3800 -6018 -3760
rect -6418 -4120 -6378 -3800
rect -6058 -4120 -6018 -3800
rect -6418 -4160 -6018 -4120
rect -5406 -3800 -5006 -3760
rect -5406 -4120 -5366 -3800
rect -5046 -4120 -5006 -3800
rect -5406 -4160 -5006 -4120
rect -4394 -3800 -3994 -3760
rect -4394 -4120 -4354 -3800
rect -4034 -4120 -3994 -3800
rect -4394 -4160 -3994 -4120
rect -3382 -3800 -2982 -3760
rect -3382 -4120 -3342 -3800
rect -3022 -4120 -2982 -3800
rect -3382 -4160 -2982 -4120
rect -2370 -3800 -1970 -3760
rect -2370 -4120 -2330 -3800
rect -2010 -4120 -1970 -3800
rect -2370 -4160 -1970 -4120
rect -1358 -3800 -958 -3760
rect -1358 -4120 -1318 -3800
rect -998 -4120 -958 -3800
rect -1358 -4160 -958 -4120
rect -346 -3800 54 -3760
rect -346 -4120 -306 -3800
rect 14 -4120 54 -3800
rect -346 -4160 54 -4120
rect 666 -3800 1066 -3760
rect 666 -4120 706 -3800
rect 1026 -4120 1066 -3800
rect 666 -4160 1066 -4120
rect 1678 -3800 2078 -3760
rect 1678 -4120 1718 -3800
rect 2038 -4120 2078 -3800
rect 1678 -4160 2078 -4120
rect 2690 -3800 3090 -3760
rect 2690 -4120 2730 -3800
rect 3050 -4120 3090 -3800
rect 2690 -4160 3090 -4120
rect 3702 -3800 4102 -3760
rect 3702 -4120 3742 -3800
rect 4062 -4120 4102 -3800
rect 3702 -4160 4102 -4120
rect 4714 -3800 5114 -3760
rect 4714 -4120 4754 -3800
rect 5074 -4120 5114 -3800
rect 4714 -4160 5114 -4120
rect 5726 -3800 6126 -3760
rect 5726 -4120 5766 -3800
rect 6086 -4120 6126 -3800
rect 5726 -4160 6126 -4120
rect 6738 -3800 7138 -3760
rect 6738 -4120 6778 -3800
rect 7098 -4120 7138 -3800
rect 6738 -4160 7138 -4120
rect -7430 -4520 -7030 -4480
rect -7430 -4840 -7390 -4520
rect -7070 -4840 -7030 -4520
rect -7430 -4880 -7030 -4840
rect -6418 -4520 -6018 -4480
rect -6418 -4840 -6378 -4520
rect -6058 -4840 -6018 -4520
rect -6418 -4880 -6018 -4840
rect -5406 -4520 -5006 -4480
rect -5406 -4840 -5366 -4520
rect -5046 -4840 -5006 -4520
rect -5406 -4880 -5006 -4840
rect -4394 -4520 -3994 -4480
rect -4394 -4840 -4354 -4520
rect -4034 -4840 -3994 -4520
rect -4394 -4880 -3994 -4840
rect -3382 -4520 -2982 -4480
rect -3382 -4840 -3342 -4520
rect -3022 -4840 -2982 -4520
rect -3382 -4880 -2982 -4840
rect -2370 -4520 -1970 -4480
rect -2370 -4840 -2330 -4520
rect -2010 -4840 -1970 -4520
rect -2370 -4880 -1970 -4840
rect -1358 -4520 -958 -4480
rect -1358 -4840 -1318 -4520
rect -998 -4840 -958 -4520
rect -1358 -4880 -958 -4840
rect -346 -4520 54 -4480
rect -346 -4840 -306 -4520
rect 14 -4840 54 -4520
rect -346 -4880 54 -4840
rect 666 -4520 1066 -4480
rect 666 -4840 706 -4520
rect 1026 -4840 1066 -4520
rect 666 -4880 1066 -4840
rect 1678 -4520 2078 -4480
rect 1678 -4840 1718 -4520
rect 2038 -4840 2078 -4520
rect 1678 -4880 2078 -4840
rect 2690 -4520 3090 -4480
rect 2690 -4840 2730 -4520
rect 3050 -4840 3090 -4520
rect 2690 -4880 3090 -4840
rect 3702 -4520 4102 -4480
rect 3702 -4840 3742 -4520
rect 4062 -4840 4102 -4520
rect 3702 -4880 4102 -4840
rect 4714 -4520 5114 -4480
rect 4714 -4840 4754 -4520
rect 5074 -4840 5114 -4520
rect 4714 -4880 5114 -4840
rect 5726 -4520 6126 -4480
rect 5726 -4840 5766 -4520
rect 6086 -4840 6126 -4520
rect 5726 -4880 6126 -4840
rect 6738 -4520 7138 -4480
rect 6738 -4840 6778 -4520
rect 7098 -4840 7138 -4520
rect 6738 -4880 7138 -4840
rect -7430 -5240 -7030 -5200
rect -7430 -5560 -7390 -5240
rect -7070 -5560 -7030 -5240
rect -7430 -5600 -7030 -5560
rect -6418 -5240 -6018 -5200
rect -6418 -5560 -6378 -5240
rect -6058 -5560 -6018 -5240
rect -6418 -5600 -6018 -5560
rect -5406 -5240 -5006 -5200
rect -5406 -5560 -5366 -5240
rect -5046 -5560 -5006 -5240
rect -5406 -5600 -5006 -5560
rect -4394 -5240 -3994 -5200
rect -4394 -5560 -4354 -5240
rect -4034 -5560 -3994 -5240
rect -4394 -5600 -3994 -5560
rect -3382 -5240 -2982 -5200
rect -3382 -5560 -3342 -5240
rect -3022 -5560 -2982 -5240
rect -3382 -5600 -2982 -5560
rect -2370 -5240 -1970 -5200
rect -2370 -5560 -2330 -5240
rect -2010 -5560 -1970 -5240
rect -2370 -5600 -1970 -5560
rect -1358 -5240 -958 -5200
rect -1358 -5560 -1318 -5240
rect -998 -5560 -958 -5240
rect -1358 -5600 -958 -5560
rect -346 -5240 54 -5200
rect -346 -5560 -306 -5240
rect 14 -5560 54 -5240
rect -346 -5600 54 -5560
rect 666 -5240 1066 -5200
rect 666 -5560 706 -5240
rect 1026 -5560 1066 -5240
rect 666 -5600 1066 -5560
rect 1678 -5240 2078 -5200
rect 1678 -5560 1718 -5240
rect 2038 -5560 2078 -5240
rect 1678 -5600 2078 -5560
rect 2690 -5240 3090 -5200
rect 2690 -5560 2730 -5240
rect 3050 -5560 3090 -5240
rect 2690 -5600 3090 -5560
rect 3702 -5240 4102 -5200
rect 3702 -5560 3742 -5240
rect 4062 -5560 4102 -5240
rect 3702 -5600 4102 -5560
rect 4714 -5240 5114 -5200
rect 4714 -5560 4754 -5240
rect 5074 -5560 5114 -5240
rect 4714 -5600 5114 -5560
rect 5726 -5240 6126 -5200
rect 5726 -5560 5766 -5240
rect 6086 -5560 6126 -5240
rect 5726 -5600 6126 -5560
rect 6738 -5240 7138 -5200
rect 6738 -5560 6778 -5240
rect 7098 -5560 7138 -5240
rect 6738 -5600 7138 -5560
rect -7430 -5960 -7030 -5920
rect -7430 -6280 -7390 -5960
rect -7070 -6280 -7030 -5960
rect -7430 -6320 -7030 -6280
rect -6418 -5960 -6018 -5920
rect -6418 -6280 -6378 -5960
rect -6058 -6280 -6018 -5960
rect -6418 -6320 -6018 -6280
rect -5406 -5960 -5006 -5920
rect -5406 -6280 -5366 -5960
rect -5046 -6280 -5006 -5960
rect -5406 -6320 -5006 -6280
rect -4394 -5960 -3994 -5920
rect -4394 -6280 -4354 -5960
rect -4034 -6280 -3994 -5960
rect -4394 -6320 -3994 -6280
rect -3382 -5960 -2982 -5920
rect -3382 -6280 -3342 -5960
rect -3022 -6280 -2982 -5960
rect -3382 -6320 -2982 -6280
rect -2370 -5960 -1970 -5920
rect -2370 -6280 -2330 -5960
rect -2010 -6280 -1970 -5960
rect -2370 -6320 -1970 -6280
rect -1358 -5960 -958 -5920
rect -1358 -6280 -1318 -5960
rect -998 -6280 -958 -5960
rect -1358 -6320 -958 -6280
rect -346 -5960 54 -5920
rect -346 -6280 -306 -5960
rect 14 -6280 54 -5960
rect -346 -6320 54 -6280
rect 666 -5960 1066 -5920
rect 666 -6280 706 -5960
rect 1026 -6280 1066 -5960
rect 666 -6320 1066 -6280
rect 1678 -5960 2078 -5920
rect 1678 -6280 1718 -5960
rect 2038 -6280 2078 -5960
rect 1678 -6320 2078 -6280
rect 2690 -5960 3090 -5920
rect 2690 -6280 2730 -5960
rect 3050 -6280 3090 -5960
rect 2690 -6320 3090 -6280
rect 3702 -5960 4102 -5920
rect 3702 -6280 3742 -5960
rect 4062 -6280 4102 -5960
rect 3702 -6320 4102 -6280
rect 4714 -5960 5114 -5920
rect 4714 -6280 4754 -5960
rect 5074 -6280 5114 -5960
rect 4714 -6320 5114 -6280
rect 5726 -5960 6126 -5920
rect 5726 -6280 5766 -5960
rect 6086 -6280 6126 -5960
rect 5726 -6320 6126 -6280
rect 6738 -5960 7138 -5920
rect 6738 -6280 6778 -5960
rect 7098 -6280 7138 -5960
rect 6738 -6320 7138 -6280
rect -7430 -6680 -7030 -6640
rect -7430 -7000 -7390 -6680
rect -7070 -7000 -7030 -6680
rect -7430 -7040 -7030 -7000
rect -6418 -6680 -6018 -6640
rect -6418 -7000 -6378 -6680
rect -6058 -7000 -6018 -6680
rect -6418 -7040 -6018 -7000
rect -5406 -6680 -5006 -6640
rect -5406 -7000 -5366 -6680
rect -5046 -7000 -5006 -6680
rect -5406 -7040 -5006 -7000
rect -4394 -6680 -3994 -6640
rect -4394 -7000 -4354 -6680
rect -4034 -7000 -3994 -6680
rect -4394 -7040 -3994 -7000
rect -3382 -6680 -2982 -6640
rect -3382 -7000 -3342 -6680
rect -3022 -7000 -2982 -6680
rect -3382 -7040 -2982 -7000
rect -2370 -6680 -1970 -6640
rect -2370 -7000 -2330 -6680
rect -2010 -7000 -1970 -6680
rect -2370 -7040 -1970 -7000
rect -1358 -6680 -958 -6640
rect -1358 -7000 -1318 -6680
rect -998 -7000 -958 -6680
rect -1358 -7040 -958 -7000
rect -346 -6680 54 -6640
rect -346 -7000 -306 -6680
rect 14 -7000 54 -6680
rect -346 -7040 54 -7000
rect 666 -6680 1066 -6640
rect 666 -7000 706 -6680
rect 1026 -7000 1066 -6680
rect 666 -7040 1066 -7000
rect 1678 -6680 2078 -6640
rect 1678 -7000 1718 -6680
rect 2038 -7000 2078 -6680
rect 1678 -7040 2078 -7000
rect 2690 -6680 3090 -6640
rect 2690 -7000 2730 -6680
rect 3050 -7000 3090 -6680
rect 2690 -7040 3090 -7000
rect 3702 -6680 4102 -6640
rect 3702 -7000 3742 -6680
rect 4062 -7000 4102 -6680
rect 3702 -7040 4102 -7000
rect 4714 -6680 5114 -6640
rect 4714 -7000 4754 -6680
rect 5074 -7000 5114 -6680
rect 4714 -7040 5114 -7000
rect 5726 -6680 6126 -6640
rect 5726 -7000 5766 -6680
rect 6086 -7000 6126 -6680
rect 5726 -7040 6126 -7000
rect 6738 -6680 7138 -6640
rect 6738 -7000 6778 -6680
rect 7098 -7000 7138 -6680
rect 6738 -7040 7138 -7000
rect -7430 -7400 -7030 -7360
rect -7430 -7720 -7390 -7400
rect -7070 -7720 -7030 -7400
rect -7430 -7760 -7030 -7720
rect -6418 -7400 -6018 -7360
rect -6418 -7720 -6378 -7400
rect -6058 -7720 -6018 -7400
rect -6418 -7760 -6018 -7720
rect -5406 -7400 -5006 -7360
rect -5406 -7720 -5366 -7400
rect -5046 -7720 -5006 -7400
rect -5406 -7760 -5006 -7720
rect -4394 -7400 -3994 -7360
rect -4394 -7720 -4354 -7400
rect -4034 -7720 -3994 -7400
rect -4394 -7760 -3994 -7720
rect -3382 -7400 -2982 -7360
rect -3382 -7720 -3342 -7400
rect -3022 -7720 -2982 -7400
rect -3382 -7760 -2982 -7720
rect -2370 -7400 -1970 -7360
rect -2370 -7720 -2330 -7400
rect -2010 -7720 -1970 -7400
rect -2370 -7760 -1970 -7720
rect -1358 -7400 -958 -7360
rect -1358 -7720 -1318 -7400
rect -998 -7720 -958 -7400
rect -1358 -7760 -958 -7720
rect -346 -7400 54 -7360
rect -346 -7720 -306 -7400
rect 14 -7720 54 -7400
rect -346 -7760 54 -7720
rect 666 -7400 1066 -7360
rect 666 -7720 706 -7400
rect 1026 -7720 1066 -7400
rect 666 -7760 1066 -7720
rect 1678 -7400 2078 -7360
rect 1678 -7720 1718 -7400
rect 2038 -7720 2078 -7400
rect 1678 -7760 2078 -7720
rect 2690 -7400 3090 -7360
rect 2690 -7720 2730 -7400
rect 3050 -7720 3090 -7400
rect 2690 -7760 3090 -7720
rect 3702 -7400 4102 -7360
rect 3702 -7720 3742 -7400
rect 4062 -7720 4102 -7400
rect 3702 -7760 4102 -7720
rect 4714 -7400 5114 -7360
rect 4714 -7720 4754 -7400
rect 5074 -7720 5114 -7400
rect 4714 -7760 5114 -7720
rect 5726 -7400 6126 -7360
rect 5726 -7720 5766 -7400
rect 6086 -7720 6126 -7400
rect 5726 -7760 6126 -7720
rect 6738 -7400 7138 -7360
rect 6738 -7720 6778 -7400
rect 7098 -7720 7138 -7400
rect 6738 -7760 7138 -7720
rect -7430 -8120 -7030 -8080
rect -7430 -8440 -7390 -8120
rect -7070 -8440 -7030 -8120
rect -7430 -8480 -7030 -8440
rect -6418 -8120 -6018 -8080
rect -6418 -8440 -6378 -8120
rect -6058 -8440 -6018 -8120
rect -6418 -8480 -6018 -8440
rect -5406 -8120 -5006 -8080
rect -5406 -8440 -5366 -8120
rect -5046 -8440 -5006 -8120
rect -5406 -8480 -5006 -8440
rect -4394 -8120 -3994 -8080
rect -4394 -8440 -4354 -8120
rect -4034 -8440 -3994 -8120
rect -4394 -8480 -3994 -8440
rect -3382 -8120 -2982 -8080
rect -3382 -8440 -3342 -8120
rect -3022 -8440 -2982 -8120
rect -3382 -8480 -2982 -8440
rect -2370 -8120 -1970 -8080
rect -2370 -8440 -2330 -8120
rect -2010 -8440 -1970 -8120
rect -2370 -8480 -1970 -8440
rect -1358 -8120 -958 -8080
rect -1358 -8440 -1318 -8120
rect -998 -8440 -958 -8120
rect -1358 -8480 -958 -8440
rect -346 -8120 54 -8080
rect -346 -8440 -306 -8120
rect 14 -8440 54 -8120
rect -346 -8480 54 -8440
rect 666 -8120 1066 -8080
rect 666 -8440 706 -8120
rect 1026 -8440 1066 -8120
rect 666 -8480 1066 -8440
rect 1678 -8120 2078 -8080
rect 1678 -8440 1718 -8120
rect 2038 -8440 2078 -8120
rect 1678 -8480 2078 -8440
rect 2690 -8120 3090 -8080
rect 2690 -8440 2730 -8120
rect 3050 -8440 3090 -8120
rect 2690 -8480 3090 -8440
rect 3702 -8120 4102 -8080
rect 3702 -8440 3742 -8120
rect 4062 -8440 4102 -8120
rect 3702 -8480 4102 -8440
rect 4714 -8120 5114 -8080
rect 4714 -8440 4754 -8120
rect 5074 -8440 5114 -8120
rect 4714 -8480 5114 -8440
rect 5726 -8120 6126 -8080
rect 5726 -8440 5766 -8120
rect 6086 -8440 6126 -8120
rect 5726 -8480 6126 -8440
rect 6738 -8120 7138 -8080
rect 6738 -8440 6778 -8120
rect 7098 -8440 7138 -8120
rect 6738 -8480 7138 -8440
rect -7430 -8840 -7030 -8800
rect -7430 -9160 -7390 -8840
rect -7070 -9160 -7030 -8840
rect -7430 -9200 -7030 -9160
rect -6418 -8840 -6018 -8800
rect -6418 -9160 -6378 -8840
rect -6058 -9160 -6018 -8840
rect -6418 -9200 -6018 -9160
rect -5406 -8840 -5006 -8800
rect -5406 -9160 -5366 -8840
rect -5046 -9160 -5006 -8840
rect -5406 -9200 -5006 -9160
rect -4394 -8840 -3994 -8800
rect -4394 -9160 -4354 -8840
rect -4034 -9160 -3994 -8840
rect -4394 -9200 -3994 -9160
rect -3382 -8840 -2982 -8800
rect -3382 -9160 -3342 -8840
rect -3022 -9160 -2982 -8840
rect -3382 -9200 -2982 -9160
rect -2370 -8840 -1970 -8800
rect -2370 -9160 -2330 -8840
rect -2010 -9160 -1970 -8840
rect -2370 -9200 -1970 -9160
rect -1358 -8840 -958 -8800
rect -1358 -9160 -1318 -8840
rect -998 -9160 -958 -8840
rect -1358 -9200 -958 -9160
rect -346 -8840 54 -8800
rect -346 -9160 -306 -8840
rect 14 -9160 54 -8840
rect -346 -9200 54 -9160
rect 666 -8840 1066 -8800
rect 666 -9160 706 -8840
rect 1026 -9160 1066 -8840
rect 666 -9200 1066 -9160
rect 1678 -8840 2078 -8800
rect 1678 -9160 1718 -8840
rect 2038 -9160 2078 -8840
rect 1678 -9200 2078 -9160
rect 2690 -8840 3090 -8800
rect 2690 -9160 2730 -8840
rect 3050 -9160 3090 -8840
rect 2690 -9200 3090 -9160
rect 3702 -8840 4102 -8800
rect 3702 -9160 3742 -8840
rect 4062 -9160 4102 -8840
rect 3702 -9200 4102 -9160
rect 4714 -8840 5114 -8800
rect 4714 -9160 4754 -8840
rect 5074 -9160 5114 -8840
rect 4714 -9200 5114 -9160
rect 5726 -8840 6126 -8800
rect 5726 -9160 5766 -8840
rect 6086 -9160 6126 -8840
rect 5726 -9200 6126 -9160
rect 6738 -8840 7138 -8800
rect 6738 -9160 6778 -8840
rect 7098 -9160 7138 -8840
rect 6738 -9200 7138 -9160
rect -7430 -9560 -7030 -9520
rect -7430 -9880 -7390 -9560
rect -7070 -9880 -7030 -9560
rect -7430 -9920 -7030 -9880
rect -6418 -9560 -6018 -9520
rect -6418 -9880 -6378 -9560
rect -6058 -9880 -6018 -9560
rect -6418 -9920 -6018 -9880
rect -5406 -9560 -5006 -9520
rect -5406 -9880 -5366 -9560
rect -5046 -9880 -5006 -9560
rect -5406 -9920 -5006 -9880
rect -4394 -9560 -3994 -9520
rect -4394 -9880 -4354 -9560
rect -4034 -9880 -3994 -9560
rect -4394 -9920 -3994 -9880
rect -3382 -9560 -2982 -9520
rect -3382 -9880 -3342 -9560
rect -3022 -9880 -2982 -9560
rect -3382 -9920 -2982 -9880
rect -2370 -9560 -1970 -9520
rect -2370 -9880 -2330 -9560
rect -2010 -9880 -1970 -9560
rect -2370 -9920 -1970 -9880
rect -1358 -9560 -958 -9520
rect -1358 -9880 -1318 -9560
rect -998 -9880 -958 -9560
rect -1358 -9920 -958 -9880
rect -346 -9560 54 -9520
rect -346 -9880 -306 -9560
rect 14 -9880 54 -9560
rect -346 -9920 54 -9880
rect 666 -9560 1066 -9520
rect 666 -9880 706 -9560
rect 1026 -9880 1066 -9560
rect 666 -9920 1066 -9880
rect 1678 -9560 2078 -9520
rect 1678 -9880 1718 -9560
rect 2038 -9880 2078 -9560
rect 1678 -9920 2078 -9880
rect 2690 -9560 3090 -9520
rect 2690 -9880 2730 -9560
rect 3050 -9880 3090 -9560
rect 2690 -9920 3090 -9880
rect 3702 -9560 4102 -9520
rect 3702 -9880 3742 -9560
rect 4062 -9880 4102 -9560
rect 3702 -9920 4102 -9880
rect 4714 -9560 5114 -9520
rect 4714 -9880 4754 -9560
rect 5074 -9880 5114 -9560
rect 4714 -9920 5114 -9880
rect 5726 -9560 6126 -9520
rect 5726 -9880 5766 -9560
rect 6086 -9880 6126 -9560
rect 5726 -9920 6126 -9880
rect 6738 -9560 7138 -9520
rect 6738 -9880 6778 -9560
rect 7098 -9880 7138 -9560
rect 6738 -9920 7138 -9880
rect -7430 -10280 -7030 -10240
rect -7430 -10600 -7390 -10280
rect -7070 -10600 -7030 -10280
rect -7430 -10640 -7030 -10600
rect -6418 -10280 -6018 -10240
rect -6418 -10600 -6378 -10280
rect -6058 -10600 -6018 -10280
rect -6418 -10640 -6018 -10600
rect -5406 -10280 -5006 -10240
rect -5406 -10600 -5366 -10280
rect -5046 -10600 -5006 -10280
rect -5406 -10640 -5006 -10600
rect -4394 -10280 -3994 -10240
rect -4394 -10600 -4354 -10280
rect -4034 -10600 -3994 -10280
rect -4394 -10640 -3994 -10600
rect -3382 -10280 -2982 -10240
rect -3382 -10600 -3342 -10280
rect -3022 -10600 -2982 -10280
rect -3382 -10640 -2982 -10600
rect -2370 -10280 -1970 -10240
rect -2370 -10600 -2330 -10280
rect -2010 -10600 -1970 -10280
rect -2370 -10640 -1970 -10600
rect -1358 -10280 -958 -10240
rect -1358 -10600 -1318 -10280
rect -998 -10600 -958 -10280
rect -1358 -10640 -958 -10600
rect -346 -10280 54 -10240
rect -346 -10600 -306 -10280
rect 14 -10600 54 -10280
rect -346 -10640 54 -10600
rect 666 -10280 1066 -10240
rect 666 -10600 706 -10280
rect 1026 -10600 1066 -10280
rect 666 -10640 1066 -10600
rect 1678 -10280 2078 -10240
rect 1678 -10600 1718 -10280
rect 2038 -10600 2078 -10280
rect 1678 -10640 2078 -10600
rect 2690 -10280 3090 -10240
rect 2690 -10600 2730 -10280
rect 3050 -10600 3090 -10280
rect 2690 -10640 3090 -10600
rect 3702 -10280 4102 -10240
rect 3702 -10600 3742 -10280
rect 4062 -10600 4102 -10280
rect 3702 -10640 4102 -10600
rect 4714 -10280 5114 -10240
rect 4714 -10600 4754 -10280
rect 5074 -10600 5114 -10280
rect 4714 -10640 5114 -10600
rect 5726 -10280 6126 -10240
rect 5726 -10600 5766 -10280
rect 6086 -10600 6126 -10280
rect 5726 -10640 6126 -10600
rect 6738 -10280 7138 -10240
rect 6738 -10600 6778 -10280
rect 7098 -10600 7138 -10280
rect 6738 -10640 7138 -10600
rect -7430 -11000 -7030 -10960
rect -7430 -11320 -7390 -11000
rect -7070 -11320 -7030 -11000
rect -7430 -11360 -7030 -11320
rect -6418 -11000 -6018 -10960
rect -6418 -11320 -6378 -11000
rect -6058 -11320 -6018 -11000
rect -6418 -11360 -6018 -11320
rect -5406 -11000 -5006 -10960
rect -5406 -11320 -5366 -11000
rect -5046 -11320 -5006 -11000
rect -5406 -11360 -5006 -11320
rect -4394 -11000 -3994 -10960
rect -4394 -11320 -4354 -11000
rect -4034 -11320 -3994 -11000
rect -4394 -11360 -3994 -11320
rect -3382 -11000 -2982 -10960
rect -3382 -11320 -3342 -11000
rect -3022 -11320 -2982 -11000
rect -3382 -11360 -2982 -11320
rect -2370 -11000 -1970 -10960
rect -2370 -11320 -2330 -11000
rect -2010 -11320 -1970 -11000
rect -2370 -11360 -1970 -11320
rect -1358 -11000 -958 -10960
rect -1358 -11320 -1318 -11000
rect -998 -11320 -958 -11000
rect -1358 -11360 -958 -11320
rect -346 -11000 54 -10960
rect -346 -11320 -306 -11000
rect 14 -11320 54 -11000
rect -346 -11360 54 -11320
rect 666 -11000 1066 -10960
rect 666 -11320 706 -11000
rect 1026 -11320 1066 -11000
rect 666 -11360 1066 -11320
rect 1678 -11000 2078 -10960
rect 1678 -11320 1718 -11000
rect 2038 -11320 2078 -11000
rect 1678 -11360 2078 -11320
rect 2690 -11000 3090 -10960
rect 2690 -11320 2730 -11000
rect 3050 -11320 3090 -11000
rect 2690 -11360 3090 -11320
rect 3702 -11000 4102 -10960
rect 3702 -11320 3742 -11000
rect 4062 -11320 4102 -11000
rect 3702 -11360 4102 -11320
rect 4714 -11000 5114 -10960
rect 4714 -11320 4754 -11000
rect 5074 -11320 5114 -11000
rect 4714 -11360 5114 -11320
rect 5726 -11000 6126 -10960
rect 5726 -11320 5766 -11000
rect 6086 -11320 6126 -11000
rect 5726 -11360 6126 -11320
rect 6738 -11000 7138 -10960
rect 6738 -11320 6778 -11000
rect 7098 -11320 7138 -11000
rect 6738 -11360 7138 -11320
<< mimcapcontact >>
rect -7390 11000 -7070 11320
rect -6378 11000 -6058 11320
rect -5366 11000 -5046 11320
rect -4354 11000 -4034 11320
rect -3342 11000 -3022 11320
rect -2330 11000 -2010 11320
rect -1318 11000 -998 11320
rect -306 11000 14 11320
rect 706 11000 1026 11320
rect 1718 11000 2038 11320
rect 2730 11000 3050 11320
rect 3742 11000 4062 11320
rect 4754 11000 5074 11320
rect 5766 11000 6086 11320
rect 6778 11000 7098 11320
rect -7390 10280 -7070 10600
rect -6378 10280 -6058 10600
rect -5366 10280 -5046 10600
rect -4354 10280 -4034 10600
rect -3342 10280 -3022 10600
rect -2330 10280 -2010 10600
rect -1318 10280 -998 10600
rect -306 10280 14 10600
rect 706 10280 1026 10600
rect 1718 10280 2038 10600
rect 2730 10280 3050 10600
rect 3742 10280 4062 10600
rect 4754 10280 5074 10600
rect 5766 10280 6086 10600
rect 6778 10280 7098 10600
rect -7390 9560 -7070 9880
rect -6378 9560 -6058 9880
rect -5366 9560 -5046 9880
rect -4354 9560 -4034 9880
rect -3342 9560 -3022 9880
rect -2330 9560 -2010 9880
rect -1318 9560 -998 9880
rect -306 9560 14 9880
rect 706 9560 1026 9880
rect 1718 9560 2038 9880
rect 2730 9560 3050 9880
rect 3742 9560 4062 9880
rect 4754 9560 5074 9880
rect 5766 9560 6086 9880
rect 6778 9560 7098 9880
rect -7390 8840 -7070 9160
rect -6378 8840 -6058 9160
rect -5366 8840 -5046 9160
rect -4354 8840 -4034 9160
rect -3342 8840 -3022 9160
rect -2330 8840 -2010 9160
rect -1318 8840 -998 9160
rect -306 8840 14 9160
rect 706 8840 1026 9160
rect 1718 8840 2038 9160
rect 2730 8840 3050 9160
rect 3742 8840 4062 9160
rect 4754 8840 5074 9160
rect 5766 8840 6086 9160
rect 6778 8840 7098 9160
rect -7390 8120 -7070 8440
rect -6378 8120 -6058 8440
rect -5366 8120 -5046 8440
rect -4354 8120 -4034 8440
rect -3342 8120 -3022 8440
rect -2330 8120 -2010 8440
rect -1318 8120 -998 8440
rect -306 8120 14 8440
rect 706 8120 1026 8440
rect 1718 8120 2038 8440
rect 2730 8120 3050 8440
rect 3742 8120 4062 8440
rect 4754 8120 5074 8440
rect 5766 8120 6086 8440
rect 6778 8120 7098 8440
rect -7390 7400 -7070 7720
rect -6378 7400 -6058 7720
rect -5366 7400 -5046 7720
rect -4354 7400 -4034 7720
rect -3342 7400 -3022 7720
rect -2330 7400 -2010 7720
rect -1318 7400 -998 7720
rect -306 7400 14 7720
rect 706 7400 1026 7720
rect 1718 7400 2038 7720
rect 2730 7400 3050 7720
rect 3742 7400 4062 7720
rect 4754 7400 5074 7720
rect 5766 7400 6086 7720
rect 6778 7400 7098 7720
rect -7390 6680 -7070 7000
rect -6378 6680 -6058 7000
rect -5366 6680 -5046 7000
rect -4354 6680 -4034 7000
rect -3342 6680 -3022 7000
rect -2330 6680 -2010 7000
rect -1318 6680 -998 7000
rect -306 6680 14 7000
rect 706 6680 1026 7000
rect 1718 6680 2038 7000
rect 2730 6680 3050 7000
rect 3742 6680 4062 7000
rect 4754 6680 5074 7000
rect 5766 6680 6086 7000
rect 6778 6680 7098 7000
rect -7390 5960 -7070 6280
rect -6378 5960 -6058 6280
rect -5366 5960 -5046 6280
rect -4354 5960 -4034 6280
rect -3342 5960 -3022 6280
rect -2330 5960 -2010 6280
rect -1318 5960 -998 6280
rect -306 5960 14 6280
rect 706 5960 1026 6280
rect 1718 5960 2038 6280
rect 2730 5960 3050 6280
rect 3742 5960 4062 6280
rect 4754 5960 5074 6280
rect 5766 5960 6086 6280
rect 6778 5960 7098 6280
rect -7390 5240 -7070 5560
rect -6378 5240 -6058 5560
rect -5366 5240 -5046 5560
rect -4354 5240 -4034 5560
rect -3342 5240 -3022 5560
rect -2330 5240 -2010 5560
rect -1318 5240 -998 5560
rect -306 5240 14 5560
rect 706 5240 1026 5560
rect 1718 5240 2038 5560
rect 2730 5240 3050 5560
rect 3742 5240 4062 5560
rect 4754 5240 5074 5560
rect 5766 5240 6086 5560
rect 6778 5240 7098 5560
rect -7390 4520 -7070 4840
rect -6378 4520 -6058 4840
rect -5366 4520 -5046 4840
rect -4354 4520 -4034 4840
rect -3342 4520 -3022 4840
rect -2330 4520 -2010 4840
rect -1318 4520 -998 4840
rect -306 4520 14 4840
rect 706 4520 1026 4840
rect 1718 4520 2038 4840
rect 2730 4520 3050 4840
rect 3742 4520 4062 4840
rect 4754 4520 5074 4840
rect 5766 4520 6086 4840
rect 6778 4520 7098 4840
rect -7390 3800 -7070 4120
rect -6378 3800 -6058 4120
rect -5366 3800 -5046 4120
rect -4354 3800 -4034 4120
rect -3342 3800 -3022 4120
rect -2330 3800 -2010 4120
rect -1318 3800 -998 4120
rect -306 3800 14 4120
rect 706 3800 1026 4120
rect 1718 3800 2038 4120
rect 2730 3800 3050 4120
rect 3742 3800 4062 4120
rect 4754 3800 5074 4120
rect 5766 3800 6086 4120
rect 6778 3800 7098 4120
rect -7390 3080 -7070 3400
rect -6378 3080 -6058 3400
rect -5366 3080 -5046 3400
rect -4354 3080 -4034 3400
rect -3342 3080 -3022 3400
rect -2330 3080 -2010 3400
rect -1318 3080 -998 3400
rect -306 3080 14 3400
rect 706 3080 1026 3400
rect 1718 3080 2038 3400
rect 2730 3080 3050 3400
rect 3742 3080 4062 3400
rect 4754 3080 5074 3400
rect 5766 3080 6086 3400
rect 6778 3080 7098 3400
rect -7390 2360 -7070 2680
rect -6378 2360 -6058 2680
rect -5366 2360 -5046 2680
rect -4354 2360 -4034 2680
rect -3342 2360 -3022 2680
rect -2330 2360 -2010 2680
rect -1318 2360 -998 2680
rect -306 2360 14 2680
rect 706 2360 1026 2680
rect 1718 2360 2038 2680
rect 2730 2360 3050 2680
rect 3742 2360 4062 2680
rect 4754 2360 5074 2680
rect 5766 2360 6086 2680
rect 6778 2360 7098 2680
rect -7390 1640 -7070 1960
rect -6378 1640 -6058 1960
rect -5366 1640 -5046 1960
rect -4354 1640 -4034 1960
rect -3342 1640 -3022 1960
rect -2330 1640 -2010 1960
rect -1318 1640 -998 1960
rect -306 1640 14 1960
rect 706 1640 1026 1960
rect 1718 1640 2038 1960
rect 2730 1640 3050 1960
rect 3742 1640 4062 1960
rect 4754 1640 5074 1960
rect 5766 1640 6086 1960
rect 6778 1640 7098 1960
rect -7390 920 -7070 1240
rect -6378 920 -6058 1240
rect -5366 920 -5046 1240
rect -4354 920 -4034 1240
rect -3342 920 -3022 1240
rect -2330 920 -2010 1240
rect -1318 920 -998 1240
rect -306 920 14 1240
rect 706 920 1026 1240
rect 1718 920 2038 1240
rect 2730 920 3050 1240
rect 3742 920 4062 1240
rect 4754 920 5074 1240
rect 5766 920 6086 1240
rect 6778 920 7098 1240
rect -7390 200 -7070 520
rect -6378 200 -6058 520
rect -5366 200 -5046 520
rect -4354 200 -4034 520
rect -3342 200 -3022 520
rect -2330 200 -2010 520
rect -1318 200 -998 520
rect -306 200 14 520
rect 706 200 1026 520
rect 1718 200 2038 520
rect 2730 200 3050 520
rect 3742 200 4062 520
rect 4754 200 5074 520
rect 5766 200 6086 520
rect 6778 200 7098 520
rect -7390 -520 -7070 -200
rect -6378 -520 -6058 -200
rect -5366 -520 -5046 -200
rect -4354 -520 -4034 -200
rect -3342 -520 -3022 -200
rect -2330 -520 -2010 -200
rect -1318 -520 -998 -200
rect -306 -520 14 -200
rect 706 -520 1026 -200
rect 1718 -520 2038 -200
rect 2730 -520 3050 -200
rect 3742 -520 4062 -200
rect 4754 -520 5074 -200
rect 5766 -520 6086 -200
rect 6778 -520 7098 -200
rect -7390 -1240 -7070 -920
rect -6378 -1240 -6058 -920
rect -5366 -1240 -5046 -920
rect -4354 -1240 -4034 -920
rect -3342 -1240 -3022 -920
rect -2330 -1240 -2010 -920
rect -1318 -1240 -998 -920
rect -306 -1240 14 -920
rect 706 -1240 1026 -920
rect 1718 -1240 2038 -920
rect 2730 -1240 3050 -920
rect 3742 -1240 4062 -920
rect 4754 -1240 5074 -920
rect 5766 -1240 6086 -920
rect 6778 -1240 7098 -920
rect -7390 -1960 -7070 -1640
rect -6378 -1960 -6058 -1640
rect -5366 -1960 -5046 -1640
rect -4354 -1960 -4034 -1640
rect -3342 -1960 -3022 -1640
rect -2330 -1960 -2010 -1640
rect -1318 -1960 -998 -1640
rect -306 -1960 14 -1640
rect 706 -1960 1026 -1640
rect 1718 -1960 2038 -1640
rect 2730 -1960 3050 -1640
rect 3742 -1960 4062 -1640
rect 4754 -1960 5074 -1640
rect 5766 -1960 6086 -1640
rect 6778 -1960 7098 -1640
rect -7390 -2680 -7070 -2360
rect -6378 -2680 -6058 -2360
rect -5366 -2680 -5046 -2360
rect -4354 -2680 -4034 -2360
rect -3342 -2680 -3022 -2360
rect -2330 -2680 -2010 -2360
rect -1318 -2680 -998 -2360
rect -306 -2680 14 -2360
rect 706 -2680 1026 -2360
rect 1718 -2680 2038 -2360
rect 2730 -2680 3050 -2360
rect 3742 -2680 4062 -2360
rect 4754 -2680 5074 -2360
rect 5766 -2680 6086 -2360
rect 6778 -2680 7098 -2360
rect -7390 -3400 -7070 -3080
rect -6378 -3400 -6058 -3080
rect -5366 -3400 -5046 -3080
rect -4354 -3400 -4034 -3080
rect -3342 -3400 -3022 -3080
rect -2330 -3400 -2010 -3080
rect -1318 -3400 -998 -3080
rect -306 -3400 14 -3080
rect 706 -3400 1026 -3080
rect 1718 -3400 2038 -3080
rect 2730 -3400 3050 -3080
rect 3742 -3400 4062 -3080
rect 4754 -3400 5074 -3080
rect 5766 -3400 6086 -3080
rect 6778 -3400 7098 -3080
rect -7390 -4120 -7070 -3800
rect -6378 -4120 -6058 -3800
rect -5366 -4120 -5046 -3800
rect -4354 -4120 -4034 -3800
rect -3342 -4120 -3022 -3800
rect -2330 -4120 -2010 -3800
rect -1318 -4120 -998 -3800
rect -306 -4120 14 -3800
rect 706 -4120 1026 -3800
rect 1718 -4120 2038 -3800
rect 2730 -4120 3050 -3800
rect 3742 -4120 4062 -3800
rect 4754 -4120 5074 -3800
rect 5766 -4120 6086 -3800
rect 6778 -4120 7098 -3800
rect -7390 -4840 -7070 -4520
rect -6378 -4840 -6058 -4520
rect -5366 -4840 -5046 -4520
rect -4354 -4840 -4034 -4520
rect -3342 -4840 -3022 -4520
rect -2330 -4840 -2010 -4520
rect -1318 -4840 -998 -4520
rect -306 -4840 14 -4520
rect 706 -4840 1026 -4520
rect 1718 -4840 2038 -4520
rect 2730 -4840 3050 -4520
rect 3742 -4840 4062 -4520
rect 4754 -4840 5074 -4520
rect 5766 -4840 6086 -4520
rect 6778 -4840 7098 -4520
rect -7390 -5560 -7070 -5240
rect -6378 -5560 -6058 -5240
rect -5366 -5560 -5046 -5240
rect -4354 -5560 -4034 -5240
rect -3342 -5560 -3022 -5240
rect -2330 -5560 -2010 -5240
rect -1318 -5560 -998 -5240
rect -306 -5560 14 -5240
rect 706 -5560 1026 -5240
rect 1718 -5560 2038 -5240
rect 2730 -5560 3050 -5240
rect 3742 -5560 4062 -5240
rect 4754 -5560 5074 -5240
rect 5766 -5560 6086 -5240
rect 6778 -5560 7098 -5240
rect -7390 -6280 -7070 -5960
rect -6378 -6280 -6058 -5960
rect -5366 -6280 -5046 -5960
rect -4354 -6280 -4034 -5960
rect -3342 -6280 -3022 -5960
rect -2330 -6280 -2010 -5960
rect -1318 -6280 -998 -5960
rect -306 -6280 14 -5960
rect 706 -6280 1026 -5960
rect 1718 -6280 2038 -5960
rect 2730 -6280 3050 -5960
rect 3742 -6280 4062 -5960
rect 4754 -6280 5074 -5960
rect 5766 -6280 6086 -5960
rect 6778 -6280 7098 -5960
rect -7390 -7000 -7070 -6680
rect -6378 -7000 -6058 -6680
rect -5366 -7000 -5046 -6680
rect -4354 -7000 -4034 -6680
rect -3342 -7000 -3022 -6680
rect -2330 -7000 -2010 -6680
rect -1318 -7000 -998 -6680
rect -306 -7000 14 -6680
rect 706 -7000 1026 -6680
rect 1718 -7000 2038 -6680
rect 2730 -7000 3050 -6680
rect 3742 -7000 4062 -6680
rect 4754 -7000 5074 -6680
rect 5766 -7000 6086 -6680
rect 6778 -7000 7098 -6680
rect -7390 -7720 -7070 -7400
rect -6378 -7720 -6058 -7400
rect -5366 -7720 -5046 -7400
rect -4354 -7720 -4034 -7400
rect -3342 -7720 -3022 -7400
rect -2330 -7720 -2010 -7400
rect -1318 -7720 -998 -7400
rect -306 -7720 14 -7400
rect 706 -7720 1026 -7400
rect 1718 -7720 2038 -7400
rect 2730 -7720 3050 -7400
rect 3742 -7720 4062 -7400
rect 4754 -7720 5074 -7400
rect 5766 -7720 6086 -7400
rect 6778 -7720 7098 -7400
rect -7390 -8440 -7070 -8120
rect -6378 -8440 -6058 -8120
rect -5366 -8440 -5046 -8120
rect -4354 -8440 -4034 -8120
rect -3342 -8440 -3022 -8120
rect -2330 -8440 -2010 -8120
rect -1318 -8440 -998 -8120
rect -306 -8440 14 -8120
rect 706 -8440 1026 -8120
rect 1718 -8440 2038 -8120
rect 2730 -8440 3050 -8120
rect 3742 -8440 4062 -8120
rect 4754 -8440 5074 -8120
rect 5766 -8440 6086 -8120
rect 6778 -8440 7098 -8120
rect -7390 -9160 -7070 -8840
rect -6378 -9160 -6058 -8840
rect -5366 -9160 -5046 -8840
rect -4354 -9160 -4034 -8840
rect -3342 -9160 -3022 -8840
rect -2330 -9160 -2010 -8840
rect -1318 -9160 -998 -8840
rect -306 -9160 14 -8840
rect 706 -9160 1026 -8840
rect 1718 -9160 2038 -8840
rect 2730 -9160 3050 -8840
rect 3742 -9160 4062 -8840
rect 4754 -9160 5074 -8840
rect 5766 -9160 6086 -8840
rect 6778 -9160 7098 -8840
rect -7390 -9880 -7070 -9560
rect -6378 -9880 -6058 -9560
rect -5366 -9880 -5046 -9560
rect -4354 -9880 -4034 -9560
rect -3342 -9880 -3022 -9560
rect -2330 -9880 -2010 -9560
rect -1318 -9880 -998 -9560
rect -306 -9880 14 -9560
rect 706 -9880 1026 -9560
rect 1718 -9880 2038 -9560
rect 2730 -9880 3050 -9560
rect 3742 -9880 4062 -9560
rect 4754 -9880 5074 -9560
rect 5766 -9880 6086 -9560
rect 6778 -9880 7098 -9560
rect -7390 -10600 -7070 -10280
rect -6378 -10600 -6058 -10280
rect -5366 -10600 -5046 -10280
rect -4354 -10600 -4034 -10280
rect -3342 -10600 -3022 -10280
rect -2330 -10600 -2010 -10280
rect -1318 -10600 -998 -10280
rect -306 -10600 14 -10280
rect 706 -10600 1026 -10280
rect 1718 -10600 2038 -10280
rect 2730 -10600 3050 -10280
rect 3742 -10600 4062 -10280
rect 4754 -10600 5074 -10280
rect 5766 -10600 6086 -10280
rect 6778 -10600 7098 -10280
rect -7390 -11320 -7070 -11000
rect -6378 -11320 -6058 -11000
rect -5366 -11320 -5046 -11000
rect -4354 -11320 -4034 -11000
rect -3342 -11320 -3022 -11000
rect -2330 -11320 -2010 -11000
rect -1318 -11320 -998 -11000
rect -306 -11320 14 -11000
rect 706 -11320 1026 -11000
rect 1718 -11320 2038 -11000
rect 2730 -11320 3050 -11000
rect 3742 -11320 4062 -11000
rect 4754 -11320 5074 -11000
rect 5766 -11320 6086 -11000
rect 6778 -11320 7098 -11000
<< metal4 >>
rect -7282 11321 -7178 11520
rect -6802 11372 -6698 11520
rect -7391 11320 -7069 11321
rect -7391 11000 -7390 11320
rect -7070 11000 -7069 11320
rect -7391 10999 -7069 11000
rect -7282 10601 -7178 10999
rect -6802 10948 -6782 11372
rect -6718 10948 -6698 11372
rect -6270 11321 -6166 11520
rect -5790 11372 -5686 11520
rect -6379 11320 -6057 11321
rect -6379 11000 -6378 11320
rect -6058 11000 -6057 11320
rect -6379 10999 -6057 11000
rect -6802 10652 -6698 10948
rect -7391 10600 -7069 10601
rect -7391 10280 -7390 10600
rect -7070 10280 -7069 10600
rect -7391 10279 -7069 10280
rect -7282 9881 -7178 10279
rect -6802 10228 -6782 10652
rect -6718 10228 -6698 10652
rect -6270 10601 -6166 10999
rect -5790 10948 -5770 11372
rect -5706 10948 -5686 11372
rect -5258 11321 -5154 11520
rect -4778 11372 -4674 11520
rect -5367 11320 -5045 11321
rect -5367 11000 -5366 11320
rect -5046 11000 -5045 11320
rect -5367 10999 -5045 11000
rect -5790 10652 -5686 10948
rect -6379 10600 -6057 10601
rect -6379 10280 -6378 10600
rect -6058 10280 -6057 10600
rect -6379 10279 -6057 10280
rect -6802 9932 -6698 10228
rect -7391 9880 -7069 9881
rect -7391 9560 -7390 9880
rect -7070 9560 -7069 9880
rect -7391 9559 -7069 9560
rect -7282 9161 -7178 9559
rect -6802 9508 -6782 9932
rect -6718 9508 -6698 9932
rect -6270 9881 -6166 10279
rect -5790 10228 -5770 10652
rect -5706 10228 -5686 10652
rect -5258 10601 -5154 10999
rect -4778 10948 -4758 11372
rect -4694 10948 -4674 11372
rect -4246 11321 -4142 11520
rect -3766 11372 -3662 11520
rect -4355 11320 -4033 11321
rect -4355 11000 -4354 11320
rect -4034 11000 -4033 11320
rect -4355 10999 -4033 11000
rect -4778 10652 -4674 10948
rect -5367 10600 -5045 10601
rect -5367 10280 -5366 10600
rect -5046 10280 -5045 10600
rect -5367 10279 -5045 10280
rect -5790 9932 -5686 10228
rect -6379 9880 -6057 9881
rect -6379 9560 -6378 9880
rect -6058 9560 -6057 9880
rect -6379 9559 -6057 9560
rect -6802 9212 -6698 9508
rect -7391 9160 -7069 9161
rect -7391 8840 -7390 9160
rect -7070 8840 -7069 9160
rect -7391 8839 -7069 8840
rect -7282 8441 -7178 8839
rect -6802 8788 -6782 9212
rect -6718 8788 -6698 9212
rect -6270 9161 -6166 9559
rect -5790 9508 -5770 9932
rect -5706 9508 -5686 9932
rect -5258 9881 -5154 10279
rect -4778 10228 -4758 10652
rect -4694 10228 -4674 10652
rect -4246 10601 -4142 10999
rect -3766 10948 -3746 11372
rect -3682 10948 -3662 11372
rect -3234 11321 -3130 11520
rect -2754 11372 -2650 11520
rect -3343 11320 -3021 11321
rect -3343 11000 -3342 11320
rect -3022 11000 -3021 11320
rect -3343 10999 -3021 11000
rect -3766 10652 -3662 10948
rect -4355 10600 -4033 10601
rect -4355 10280 -4354 10600
rect -4034 10280 -4033 10600
rect -4355 10279 -4033 10280
rect -4778 9932 -4674 10228
rect -5367 9880 -5045 9881
rect -5367 9560 -5366 9880
rect -5046 9560 -5045 9880
rect -5367 9559 -5045 9560
rect -5790 9212 -5686 9508
rect -6379 9160 -6057 9161
rect -6379 8840 -6378 9160
rect -6058 8840 -6057 9160
rect -6379 8839 -6057 8840
rect -6802 8492 -6698 8788
rect -7391 8440 -7069 8441
rect -7391 8120 -7390 8440
rect -7070 8120 -7069 8440
rect -7391 8119 -7069 8120
rect -7282 7721 -7178 8119
rect -6802 8068 -6782 8492
rect -6718 8068 -6698 8492
rect -6270 8441 -6166 8839
rect -5790 8788 -5770 9212
rect -5706 8788 -5686 9212
rect -5258 9161 -5154 9559
rect -4778 9508 -4758 9932
rect -4694 9508 -4674 9932
rect -4246 9881 -4142 10279
rect -3766 10228 -3746 10652
rect -3682 10228 -3662 10652
rect -3234 10601 -3130 10999
rect -2754 10948 -2734 11372
rect -2670 10948 -2650 11372
rect -2222 11321 -2118 11520
rect -1742 11372 -1638 11520
rect -2331 11320 -2009 11321
rect -2331 11000 -2330 11320
rect -2010 11000 -2009 11320
rect -2331 10999 -2009 11000
rect -2754 10652 -2650 10948
rect -3343 10600 -3021 10601
rect -3343 10280 -3342 10600
rect -3022 10280 -3021 10600
rect -3343 10279 -3021 10280
rect -3766 9932 -3662 10228
rect -4355 9880 -4033 9881
rect -4355 9560 -4354 9880
rect -4034 9560 -4033 9880
rect -4355 9559 -4033 9560
rect -4778 9212 -4674 9508
rect -5367 9160 -5045 9161
rect -5367 8840 -5366 9160
rect -5046 8840 -5045 9160
rect -5367 8839 -5045 8840
rect -5790 8492 -5686 8788
rect -6379 8440 -6057 8441
rect -6379 8120 -6378 8440
rect -6058 8120 -6057 8440
rect -6379 8119 -6057 8120
rect -6802 7772 -6698 8068
rect -7391 7720 -7069 7721
rect -7391 7400 -7390 7720
rect -7070 7400 -7069 7720
rect -7391 7399 -7069 7400
rect -7282 7001 -7178 7399
rect -6802 7348 -6782 7772
rect -6718 7348 -6698 7772
rect -6270 7721 -6166 8119
rect -5790 8068 -5770 8492
rect -5706 8068 -5686 8492
rect -5258 8441 -5154 8839
rect -4778 8788 -4758 9212
rect -4694 8788 -4674 9212
rect -4246 9161 -4142 9559
rect -3766 9508 -3746 9932
rect -3682 9508 -3662 9932
rect -3234 9881 -3130 10279
rect -2754 10228 -2734 10652
rect -2670 10228 -2650 10652
rect -2222 10601 -2118 10999
rect -1742 10948 -1722 11372
rect -1658 10948 -1638 11372
rect -1210 11321 -1106 11520
rect -730 11372 -626 11520
rect -1319 11320 -997 11321
rect -1319 11000 -1318 11320
rect -998 11000 -997 11320
rect -1319 10999 -997 11000
rect -1742 10652 -1638 10948
rect -2331 10600 -2009 10601
rect -2331 10280 -2330 10600
rect -2010 10280 -2009 10600
rect -2331 10279 -2009 10280
rect -2754 9932 -2650 10228
rect -3343 9880 -3021 9881
rect -3343 9560 -3342 9880
rect -3022 9560 -3021 9880
rect -3343 9559 -3021 9560
rect -3766 9212 -3662 9508
rect -4355 9160 -4033 9161
rect -4355 8840 -4354 9160
rect -4034 8840 -4033 9160
rect -4355 8839 -4033 8840
rect -4778 8492 -4674 8788
rect -5367 8440 -5045 8441
rect -5367 8120 -5366 8440
rect -5046 8120 -5045 8440
rect -5367 8119 -5045 8120
rect -5790 7772 -5686 8068
rect -6379 7720 -6057 7721
rect -6379 7400 -6378 7720
rect -6058 7400 -6057 7720
rect -6379 7399 -6057 7400
rect -6802 7052 -6698 7348
rect -7391 7000 -7069 7001
rect -7391 6680 -7390 7000
rect -7070 6680 -7069 7000
rect -7391 6679 -7069 6680
rect -7282 6281 -7178 6679
rect -6802 6628 -6782 7052
rect -6718 6628 -6698 7052
rect -6270 7001 -6166 7399
rect -5790 7348 -5770 7772
rect -5706 7348 -5686 7772
rect -5258 7721 -5154 8119
rect -4778 8068 -4758 8492
rect -4694 8068 -4674 8492
rect -4246 8441 -4142 8839
rect -3766 8788 -3746 9212
rect -3682 8788 -3662 9212
rect -3234 9161 -3130 9559
rect -2754 9508 -2734 9932
rect -2670 9508 -2650 9932
rect -2222 9881 -2118 10279
rect -1742 10228 -1722 10652
rect -1658 10228 -1638 10652
rect -1210 10601 -1106 10999
rect -730 10948 -710 11372
rect -646 10948 -626 11372
rect -198 11321 -94 11520
rect 282 11372 386 11520
rect -307 11320 15 11321
rect -307 11000 -306 11320
rect 14 11000 15 11320
rect -307 10999 15 11000
rect -730 10652 -626 10948
rect -1319 10600 -997 10601
rect -1319 10280 -1318 10600
rect -998 10280 -997 10600
rect -1319 10279 -997 10280
rect -1742 9932 -1638 10228
rect -2331 9880 -2009 9881
rect -2331 9560 -2330 9880
rect -2010 9560 -2009 9880
rect -2331 9559 -2009 9560
rect -2754 9212 -2650 9508
rect -3343 9160 -3021 9161
rect -3343 8840 -3342 9160
rect -3022 8840 -3021 9160
rect -3343 8839 -3021 8840
rect -3766 8492 -3662 8788
rect -4355 8440 -4033 8441
rect -4355 8120 -4354 8440
rect -4034 8120 -4033 8440
rect -4355 8119 -4033 8120
rect -4778 7772 -4674 8068
rect -5367 7720 -5045 7721
rect -5367 7400 -5366 7720
rect -5046 7400 -5045 7720
rect -5367 7399 -5045 7400
rect -5790 7052 -5686 7348
rect -6379 7000 -6057 7001
rect -6379 6680 -6378 7000
rect -6058 6680 -6057 7000
rect -6379 6679 -6057 6680
rect -6802 6332 -6698 6628
rect -7391 6280 -7069 6281
rect -7391 5960 -7390 6280
rect -7070 5960 -7069 6280
rect -7391 5959 -7069 5960
rect -7282 5561 -7178 5959
rect -6802 5908 -6782 6332
rect -6718 5908 -6698 6332
rect -6270 6281 -6166 6679
rect -5790 6628 -5770 7052
rect -5706 6628 -5686 7052
rect -5258 7001 -5154 7399
rect -4778 7348 -4758 7772
rect -4694 7348 -4674 7772
rect -4246 7721 -4142 8119
rect -3766 8068 -3746 8492
rect -3682 8068 -3662 8492
rect -3234 8441 -3130 8839
rect -2754 8788 -2734 9212
rect -2670 8788 -2650 9212
rect -2222 9161 -2118 9559
rect -1742 9508 -1722 9932
rect -1658 9508 -1638 9932
rect -1210 9881 -1106 10279
rect -730 10228 -710 10652
rect -646 10228 -626 10652
rect -198 10601 -94 10999
rect 282 10948 302 11372
rect 366 10948 386 11372
rect 814 11321 918 11520
rect 1294 11372 1398 11520
rect 705 11320 1027 11321
rect 705 11000 706 11320
rect 1026 11000 1027 11320
rect 705 10999 1027 11000
rect 282 10652 386 10948
rect -307 10600 15 10601
rect -307 10280 -306 10600
rect 14 10280 15 10600
rect -307 10279 15 10280
rect -730 9932 -626 10228
rect -1319 9880 -997 9881
rect -1319 9560 -1318 9880
rect -998 9560 -997 9880
rect -1319 9559 -997 9560
rect -1742 9212 -1638 9508
rect -2331 9160 -2009 9161
rect -2331 8840 -2330 9160
rect -2010 8840 -2009 9160
rect -2331 8839 -2009 8840
rect -2754 8492 -2650 8788
rect -3343 8440 -3021 8441
rect -3343 8120 -3342 8440
rect -3022 8120 -3021 8440
rect -3343 8119 -3021 8120
rect -3766 7772 -3662 8068
rect -4355 7720 -4033 7721
rect -4355 7400 -4354 7720
rect -4034 7400 -4033 7720
rect -4355 7399 -4033 7400
rect -4778 7052 -4674 7348
rect -5367 7000 -5045 7001
rect -5367 6680 -5366 7000
rect -5046 6680 -5045 7000
rect -5367 6679 -5045 6680
rect -5790 6332 -5686 6628
rect -6379 6280 -6057 6281
rect -6379 5960 -6378 6280
rect -6058 5960 -6057 6280
rect -6379 5959 -6057 5960
rect -6802 5612 -6698 5908
rect -7391 5560 -7069 5561
rect -7391 5240 -7390 5560
rect -7070 5240 -7069 5560
rect -7391 5239 -7069 5240
rect -7282 4841 -7178 5239
rect -6802 5188 -6782 5612
rect -6718 5188 -6698 5612
rect -6270 5561 -6166 5959
rect -5790 5908 -5770 6332
rect -5706 5908 -5686 6332
rect -5258 6281 -5154 6679
rect -4778 6628 -4758 7052
rect -4694 6628 -4674 7052
rect -4246 7001 -4142 7399
rect -3766 7348 -3746 7772
rect -3682 7348 -3662 7772
rect -3234 7721 -3130 8119
rect -2754 8068 -2734 8492
rect -2670 8068 -2650 8492
rect -2222 8441 -2118 8839
rect -1742 8788 -1722 9212
rect -1658 8788 -1638 9212
rect -1210 9161 -1106 9559
rect -730 9508 -710 9932
rect -646 9508 -626 9932
rect -198 9881 -94 10279
rect 282 10228 302 10652
rect 366 10228 386 10652
rect 814 10601 918 10999
rect 1294 10948 1314 11372
rect 1378 10948 1398 11372
rect 1826 11321 1930 11520
rect 2306 11372 2410 11520
rect 1717 11320 2039 11321
rect 1717 11000 1718 11320
rect 2038 11000 2039 11320
rect 1717 10999 2039 11000
rect 1294 10652 1398 10948
rect 705 10600 1027 10601
rect 705 10280 706 10600
rect 1026 10280 1027 10600
rect 705 10279 1027 10280
rect 282 9932 386 10228
rect -307 9880 15 9881
rect -307 9560 -306 9880
rect 14 9560 15 9880
rect -307 9559 15 9560
rect -730 9212 -626 9508
rect -1319 9160 -997 9161
rect -1319 8840 -1318 9160
rect -998 8840 -997 9160
rect -1319 8839 -997 8840
rect -1742 8492 -1638 8788
rect -2331 8440 -2009 8441
rect -2331 8120 -2330 8440
rect -2010 8120 -2009 8440
rect -2331 8119 -2009 8120
rect -2754 7772 -2650 8068
rect -3343 7720 -3021 7721
rect -3343 7400 -3342 7720
rect -3022 7400 -3021 7720
rect -3343 7399 -3021 7400
rect -3766 7052 -3662 7348
rect -4355 7000 -4033 7001
rect -4355 6680 -4354 7000
rect -4034 6680 -4033 7000
rect -4355 6679 -4033 6680
rect -4778 6332 -4674 6628
rect -5367 6280 -5045 6281
rect -5367 5960 -5366 6280
rect -5046 5960 -5045 6280
rect -5367 5959 -5045 5960
rect -5790 5612 -5686 5908
rect -6379 5560 -6057 5561
rect -6379 5240 -6378 5560
rect -6058 5240 -6057 5560
rect -6379 5239 -6057 5240
rect -6802 4892 -6698 5188
rect -7391 4840 -7069 4841
rect -7391 4520 -7390 4840
rect -7070 4520 -7069 4840
rect -7391 4519 -7069 4520
rect -7282 4121 -7178 4519
rect -6802 4468 -6782 4892
rect -6718 4468 -6698 4892
rect -6270 4841 -6166 5239
rect -5790 5188 -5770 5612
rect -5706 5188 -5686 5612
rect -5258 5561 -5154 5959
rect -4778 5908 -4758 6332
rect -4694 5908 -4674 6332
rect -4246 6281 -4142 6679
rect -3766 6628 -3746 7052
rect -3682 6628 -3662 7052
rect -3234 7001 -3130 7399
rect -2754 7348 -2734 7772
rect -2670 7348 -2650 7772
rect -2222 7721 -2118 8119
rect -1742 8068 -1722 8492
rect -1658 8068 -1638 8492
rect -1210 8441 -1106 8839
rect -730 8788 -710 9212
rect -646 8788 -626 9212
rect -198 9161 -94 9559
rect 282 9508 302 9932
rect 366 9508 386 9932
rect 814 9881 918 10279
rect 1294 10228 1314 10652
rect 1378 10228 1398 10652
rect 1826 10601 1930 10999
rect 2306 10948 2326 11372
rect 2390 10948 2410 11372
rect 2838 11321 2942 11520
rect 3318 11372 3422 11520
rect 2729 11320 3051 11321
rect 2729 11000 2730 11320
rect 3050 11000 3051 11320
rect 2729 10999 3051 11000
rect 2306 10652 2410 10948
rect 1717 10600 2039 10601
rect 1717 10280 1718 10600
rect 2038 10280 2039 10600
rect 1717 10279 2039 10280
rect 1294 9932 1398 10228
rect 705 9880 1027 9881
rect 705 9560 706 9880
rect 1026 9560 1027 9880
rect 705 9559 1027 9560
rect 282 9212 386 9508
rect -307 9160 15 9161
rect -307 8840 -306 9160
rect 14 8840 15 9160
rect -307 8839 15 8840
rect -730 8492 -626 8788
rect -1319 8440 -997 8441
rect -1319 8120 -1318 8440
rect -998 8120 -997 8440
rect -1319 8119 -997 8120
rect -1742 7772 -1638 8068
rect -2331 7720 -2009 7721
rect -2331 7400 -2330 7720
rect -2010 7400 -2009 7720
rect -2331 7399 -2009 7400
rect -2754 7052 -2650 7348
rect -3343 7000 -3021 7001
rect -3343 6680 -3342 7000
rect -3022 6680 -3021 7000
rect -3343 6679 -3021 6680
rect -3766 6332 -3662 6628
rect -4355 6280 -4033 6281
rect -4355 5960 -4354 6280
rect -4034 5960 -4033 6280
rect -4355 5959 -4033 5960
rect -4778 5612 -4674 5908
rect -5367 5560 -5045 5561
rect -5367 5240 -5366 5560
rect -5046 5240 -5045 5560
rect -5367 5239 -5045 5240
rect -5790 4892 -5686 5188
rect -6379 4840 -6057 4841
rect -6379 4520 -6378 4840
rect -6058 4520 -6057 4840
rect -6379 4519 -6057 4520
rect -6802 4172 -6698 4468
rect -7391 4120 -7069 4121
rect -7391 3800 -7390 4120
rect -7070 3800 -7069 4120
rect -7391 3799 -7069 3800
rect -7282 3401 -7178 3799
rect -6802 3748 -6782 4172
rect -6718 3748 -6698 4172
rect -6270 4121 -6166 4519
rect -5790 4468 -5770 4892
rect -5706 4468 -5686 4892
rect -5258 4841 -5154 5239
rect -4778 5188 -4758 5612
rect -4694 5188 -4674 5612
rect -4246 5561 -4142 5959
rect -3766 5908 -3746 6332
rect -3682 5908 -3662 6332
rect -3234 6281 -3130 6679
rect -2754 6628 -2734 7052
rect -2670 6628 -2650 7052
rect -2222 7001 -2118 7399
rect -1742 7348 -1722 7772
rect -1658 7348 -1638 7772
rect -1210 7721 -1106 8119
rect -730 8068 -710 8492
rect -646 8068 -626 8492
rect -198 8441 -94 8839
rect 282 8788 302 9212
rect 366 8788 386 9212
rect 814 9161 918 9559
rect 1294 9508 1314 9932
rect 1378 9508 1398 9932
rect 1826 9881 1930 10279
rect 2306 10228 2326 10652
rect 2390 10228 2410 10652
rect 2838 10601 2942 10999
rect 3318 10948 3338 11372
rect 3402 10948 3422 11372
rect 3850 11321 3954 11520
rect 4330 11372 4434 11520
rect 3741 11320 4063 11321
rect 3741 11000 3742 11320
rect 4062 11000 4063 11320
rect 3741 10999 4063 11000
rect 3318 10652 3422 10948
rect 2729 10600 3051 10601
rect 2729 10280 2730 10600
rect 3050 10280 3051 10600
rect 2729 10279 3051 10280
rect 2306 9932 2410 10228
rect 1717 9880 2039 9881
rect 1717 9560 1718 9880
rect 2038 9560 2039 9880
rect 1717 9559 2039 9560
rect 1294 9212 1398 9508
rect 705 9160 1027 9161
rect 705 8840 706 9160
rect 1026 8840 1027 9160
rect 705 8839 1027 8840
rect 282 8492 386 8788
rect -307 8440 15 8441
rect -307 8120 -306 8440
rect 14 8120 15 8440
rect -307 8119 15 8120
rect -730 7772 -626 8068
rect -1319 7720 -997 7721
rect -1319 7400 -1318 7720
rect -998 7400 -997 7720
rect -1319 7399 -997 7400
rect -1742 7052 -1638 7348
rect -2331 7000 -2009 7001
rect -2331 6680 -2330 7000
rect -2010 6680 -2009 7000
rect -2331 6679 -2009 6680
rect -2754 6332 -2650 6628
rect -3343 6280 -3021 6281
rect -3343 5960 -3342 6280
rect -3022 5960 -3021 6280
rect -3343 5959 -3021 5960
rect -3766 5612 -3662 5908
rect -4355 5560 -4033 5561
rect -4355 5240 -4354 5560
rect -4034 5240 -4033 5560
rect -4355 5239 -4033 5240
rect -4778 4892 -4674 5188
rect -5367 4840 -5045 4841
rect -5367 4520 -5366 4840
rect -5046 4520 -5045 4840
rect -5367 4519 -5045 4520
rect -5790 4172 -5686 4468
rect -6379 4120 -6057 4121
rect -6379 3800 -6378 4120
rect -6058 3800 -6057 4120
rect -6379 3799 -6057 3800
rect -6802 3452 -6698 3748
rect -7391 3400 -7069 3401
rect -7391 3080 -7390 3400
rect -7070 3080 -7069 3400
rect -7391 3079 -7069 3080
rect -7282 2681 -7178 3079
rect -6802 3028 -6782 3452
rect -6718 3028 -6698 3452
rect -6270 3401 -6166 3799
rect -5790 3748 -5770 4172
rect -5706 3748 -5686 4172
rect -5258 4121 -5154 4519
rect -4778 4468 -4758 4892
rect -4694 4468 -4674 4892
rect -4246 4841 -4142 5239
rect -3766 5188 -3746 5612
rect -3682 5188 -3662 5612
rect -3234 5561 -3130 5959
rect -2754 5908 -2734 6332
rect -2670 5908 -2650 6332
rect -2222 6281 -2118 6679
rect -1742 6628 -1722 7052
rect -1658 6628 -1638 7052
rect -1210 7001 -1106 7399
rect -730 7348 -710 7772
rect -646 7348 -626 7772
rect -198 7721 -94 8119
rect 282 8068 302 8492
rect 366 8068 386 8492
rect 814 8441 918 8839
rect 1294 8788 1314 9212
rect 1378 8788 1398 9212
rect 1826 9161 1930 9559
rect 2306 9508 2326 9932
rect 2390 9508 2410 9932
rect 2838 9881 2942 10279
rect 3318 10228 3338 10652
rect 3402 10228 3422 10652
rect 3850 10601 3954 10999
rect 4330 10948 4350 11372
rect 4414 10948 4434 11372
rect 4862 11321 4966 11520
rect 5342 11372 5446 11520
rect 4753 11320 5075 11321
rect 4753 11000 4754 11320
rect 5074 11000 5075 11320
rect 4753 10999 5075 11000
rect 4330 10652 4434 10948
rect 3741 10600 4063 10601
rect 3741 10280 3742 10600
rect 4062 10280 4063 10600
rect 3741 10279 4063 10280
rect 3318 9932 3422 10228
rect 2729 9880 3051 9881
rect 2729 9560 2730 9880
rect 3050 9560 3051 9880
rect 2729 9559 3051 9560
rect 2306 9212 2410 9508
rect 1717 9160 2039 9161
rect 1717 8840 1718 9160
rect 2038 8840 2039 9160
rect 1717 8839 2039 8840
rect 1294 8492 1398 8788
rect 705 8440 1027 8441
rect 705 8120 706 8440
rect 1026 8120 1027 8440
rect 705 8119 1027 8120
rect 282 7772 386 8068
rect -307 7720 15 7721
rect -307 7400 -306 7720
rect 14 7400 15 7720
rect -307 7399 15 7400
rect -730 7052 -626 7348
rect -1319 7000 -997 7001
rect -1319 6680 -1318 7000
rect -998 6680 -997 7000
rect -1319 6679 -997 6680
rect -1742 6332 -1638 6628
rect -2331 6280 -2009 6281
rect -2331 5960 -2330 6280
rect -2010 5960 -2009 6280
rect -2331 5959 -2009 5960
rect -2754 5612 -2650 5908
rect -3343 5560 -3021 5561
rect -3343 5240 -3342 5560
rect -3022 5240 -3021 5560
rect -3343 5239 -3021 5240
rect -3766 4892 -3662 5188
rect -4355 4840 -4033 4841
rect -4355 4520 -4354 4840
rect -4034 4520 -4033 4840
rect -4355 4519 -4033 4520
rect -4778 4172 -4674 4468
rect -5367 4120 -5045 4121
rect -5367 3800 -5366 4120
rect -5046 3800 -5045 4120
rect -5367 3799 -5045 3800
rect -5790 3452 -5686 3748
rect -6379 3400 -6057 3401
rect -6379 3080 -6378 3400
rect -6058 3080 -6057 3400
rect -6379 3079 -6057 3080
rect -6802 2732 -6698 3028
rect -7391 2680 -7069 2681
rect -7391 2360 -7390 2680
rect -7070 2360 -7069 2680
rect -7391 2359 -7069 2360
rect -7282 1961 -7178 2359
rect -6802 2308 -6782 2732
rect -6718 2308 -6698 2732
rect -6270 2681 -6166 3079
rect -5790 3028 -5770 3452
rect -5706 3028 -5686 3452
rect -5258 3401 -5154 3799
rect -4778 3748 -4758 4172
rect -4694 3748 -4674 4172
rect -4246 4121 -4142 4519
rect -3766 4468 -3746 4892
rect -3682 4468 -3662 4892
rect -3234 4841 -3130 5239
rect -2754 5188 -2734 5612
rect -2670 5188 -2650 5612
rect -2222 5561 -2118 5959
rect -1742 5908 -1722 6332
rect -1658 5908 -1638 6332
rect -1210 6281 -1106 6679
rect -730 6628 -710 7052
rect -646 6628 -626 7052
rect -198 7001 -94 7399
rect 282 7348 302 7772
rect 366 7348 386 7772
rect 814 7721 918 8119
rect 1294 8068 1314 8492
rect 1378 8068 1398 8492
rect 1826 8441 1930 8839
rect 2306 8788 2326 9212
rect 2390 8788 2410 9212
rect 2838 9161 2942 9559
rect 3318 9508 3338 9932
rect 3402 9508 3422 9932
rect 3850 9881 3954 10279
rect 4330 10228 4350 10652
rect 4414 10228 4434 10652
rect 4862 10601 4966 10999
rect 5342 10948 5362 11372
rect 5426 10948 5446 11372
rect 5874 11321 5978 11520
rect 6354 11372 6458 11520
rect 5765 11320 6087 11321
rect 5765 11000 5766 11320
rect 6086 11000 6087 11320
rect 5765 10999 6087 11000
rect 5342 10652 5446 10948
rect 4753 10600 5075 10601
rect 4753 10280 4754 10600
rect 5074 10280 5075 10600
rect 4753 10279 5075 10280
rect 4330 9932 4434 10228
rect 3741 9880 4063 9881
rect 3741 9560 3742 9880
rect 4062 9560 4063 9880
rect 3741 9559 4063 9560
rect 3318 9212 3422 9508
rect 2729 9160 3051 9161
rect 2729 8840 2730 9160
rect 3050 8840 3051 9160
rect 2729 8839 3051 8840
rect 2306 8492 2410 8788
rect 1717 8440 2039 8441
rect 1717 8120 1718 8440
rect 2038 8120 2039 8440
rect 1717 8119 2039 8120
rect 1294 7772 1398 8068
rect 705 7720 1027 7721
rect 705 7400 706 7720
rect 1026 7400 1027 7720
rect 705 7399 1027 7400
rect 282 7052 386 7348
rect -307 7000 15 7001
rect -307 6680 -306 7000
rect 14 6680 15 7000
rect -307 6679 15 6680
rect -730 6332 -626 6628
rect -1319 6280 -997 6281
rect -1319 5960 -1318 6280
rect -998 5960 -997 6280
rect -1319 5959 -997 5960
rect -1742 5612 -1638 5908
rect -2331 5560 -2009 5561
rect -2331 5240 -2330 5560
rect -2010 5240 -2009 5560
rect -2331 5239 -2009 5240
rect -2754 4892 -2650 5188
rect -3343 4840 -3021 4841
rect -3343 4520 -3342 4840
rect -3022 4520 -3021 4840
rect -3343 4519 -3021 4520
rect -3766 4172 -3662 4468
rect -4355 4120 -4033 4121
rect -4355 3800 -4354 4120
rect -4034 3800 -4033 4120
rect -4355 3799 -4033 3800
rect -4778 3452 -4674 3748
rect -5367 3400 -5045 3401
rect -5367 3080 -5366 3400
rect -5046 3080 -5045 3400
rect -5367 3079 -5045 3080
rect -5790 2732 -5686 3028
rect -6379 2680 -6057 2681
rect -6379 2360 -6378 2680
rect -6058 2360 -6057 2680
rect -6379 2359 -6057 2360
rect -6802 2012 -6698 2308
rect -7391 1960 -7069 1961
rect -7391 1640 -7390 1960
rect -7070 1640 -7069 1960
rect -7391 1639 -7069 1640
rect -7282 1241 -7178 1639
rect -6802 1588 -6782 2012
rect -6718 1588 -6698 2012
rect -6270 1961 -6166 2359
rect -5790 2308 -5770 2732
rect -5706 2308 -5686 2732
rect -5258 2681 -5154 3079
rect -4778 3028 -4758 3452
rect -4694 3028 -4674 3452
rect -4246 3401 -4142 3799
rect -3766 3748 -3746 4172
rect -3682 3748 -3662 4172
rect -3234 4121 -3130 4519
rect -2754 4468 -2734 4892
rect -2670 4468 -2650 4892
rect -2222 4841 -2118 5239
rect -1742 5188 -1722 5612
rect -1658 5188 -1638 5612
rect -1210 5561 -1106 5959
rect -730 5908 -710 6332
rect -646 5908 -626 6332
rect -198 6281 -94 6679
rect 282 6628 302 7052
rect 366 6628 386 7052
rect 814 7001 918 7399
rect 1294 7348 1314 7772
rect 1378 7348 1398 7772
rect 1826 7721 1930 8119
rect 2306 8068 2326 8492
rect 2390 8068 2410 8492
rect 2838 8441 2942 8839
rect 3318 8788 3338 9212
rect 3402 8788 3422 9212
rect 3850 9161 3954 9559
rect 4330 9508 4350 9932
rect 4414 9508 4434 9932
rect 4862 9881 4966 10279
rect 5342 10228 5362 10652
rect 5426 10228 5446 10652
rect 5874 10601 5978 10999
rect 6354 10948 6374 11372
rect 6438 10948 6458 11372
rect 6886 11321 6990 11520
rect 7366 11372 7470 11520
rect 6777 11320 7099 11321
rect 6777 11000 6778 11320
rect 7098 11000 7099 11320
rect 6777 10999 7099 11000
rect 6354 10652 6458 10948
rect 5765 10600 6087 10601
rect 5765 10280 5766 10600
rect 6086 10280 6087 10600
rect 5765 10279 6087 10280
rect 5342 9932 5446 10228
rect 4753 9880 5075 9881
rect 4753 9560 4754 9880
rect 5074 9560 5075 9880
rect 4753 9559 5075 9560
rect 4330 9212 4434 9508
rect 3741 9160 4063 9161
rect 3741 8840 3742 9160
rect 4062 8840 4063 9160
rect 3741 8839 4063 8840
rect 3318 8492 3422 8788
rect 2729 8440 3051 8441
rect 2729 8120 2730 8440
rect 3050 8120 3051 8440
rect 2729 8119 3051 8120
rect 2306 7772 2410 8068
rect 1717 7720 2039 7721
rect 1717 7400 1718 7720
rect 2038 7400 2039 7720
rect 1717 7399 2039 7400
rect 1294 7052 1398 7348
rect 705 7000 1027 7001
rect 705 6680 706 7000
rect 1026 6680 1027 7000
rect 705 6679 1027 6680
rect 282 6332 386 6628
rect -307 6280 15 6281
rect -307 5960 -306 6280
rect 14 5960 15 6280
rect -307 5959 15 5960
rect -730 5612 -626 5908
rect -1319 5560 -997 5561
rect -1319 5240 -1318 5560
rect -998 5240 -997 5560
rect -1319 5239 -997 5240
rect -1742 4892 -1638 5188
rect -2331 4840 -2009 4841
rect -2331 4520 -2330 4840
rect -2010 4520 -2009 4840
rect -2331 4519 -2009 4520
rect -2754 4172 -2650 4468
rect -3343 4120 -3021 4121
rect -3343 3800 -3342 4120
rect -3022 3800 -3021 4120
rect -3343 3799 -3021 3800
rect -3766 3452 -3662 3748
rect -4355 3400 -4033 3401
rect -4355 3080 -4354 3400
rect -4034 3080 -4033 3400
rect -4355 3079 -4033 3080
rect -4778 2732 -4674 3028
rect -5367 2680 -5045 2681
rect -5367 2360 -5366 2680
rect -5046 2360 -5045 2680
rect -5367 2359 -5045 2360
rect -5790 2012 -5686 2308
rect -6379 1960 -6057 1961
rect -6379 1640 -6378 1960
rect -6058 1640 -6057 1960
rect -6379 1639 -6057 1640
rect -6802 1292 -6698 1588
rect -7391 1240 -7069 1241
rect -7391 920 -7390 1240
rect -7070 920 -7069 1240
rect -7391 919 -7069 920
rect -7282 521 -7178 919
rect -6802 868 -6782 1292
rect -6718 868 -6698 1292
rect -6270 1241 -6166 1639
rect -5790 1588 -5770 2012
rect -5706 1588 -5686 2012
rect -5258 1961 -5154 2359
rect -4778 2308 -4758 2732
rect -4694 2308 -4674 2732
rect -4246 2681 -4142 3079
rect -3766 3028 -3746 3452
rect -3682 3028 -3662 3452
rect -3234 3401 -3130 3799
rect -2754 3748 -2734 4172
rect -2670 3748 -2650 4172
rect -2222 4121 -2118 4519
rect -1742 4468 -1722 4892
rect -1658 4468 -1638 4892
rect -1210 4841 -1106 5239
rect -730 5188 -710 5612
rect -646 5188 -626 5612
rect -198 5561 -94 5959
rect 282 5908 302 6332
rect 366 5908 386 6332
rect 814 6281 918 6679
rect 1294 6628 1314 7052
rect 1378 6628 1398 7052
rect 1826 7001 1930 7399
rect 2306 7348 2326 7772
rect 2390 7348 2410 7772
rect 2838 7721 2942 8119
rect 3318 8068 3338 8492
rect 3402 8068 3422 8492
rect 3850 8441 3954 8839
rect 4330 8788 4350 9212
rect 4414 8788 4434 9212
rect 4862 9161 4966 9559
rect 5342 9508 5362 9932
rect 5426 9508 5446 9932
rect 5874 9881 5978 10279
rect 6354 10228 6374 10652
rect 6438 10228 6458 10652
rect 6886 10601 6990 10999
rect 7366 10948 7386 11372
rect 7450 10948 7470 11372
rect 7366 10652 7470 10948
rect 6777 10600 7099 10601
rect 6777 10280 6778 10600
rect 7098 10280 7099 10600
rect 6777 10279 7099 10280
rect 6354 9932 6458 10228
rect 5765 9880 6087 9881
rect 5765 9560 5766 9880
rect 6086 9560 6087 9880
rect 5765 9559 6087 9560
rect 5342 9212 5446 9508
rect 4753 9160 5075 9161
rect 4753 8840 4754 9160
rect 5074 8840 5075 9160
rect 4753 8839 5075 8840
rect 4330 8492 4434 8788
rect 3741 8440 4063 8441
rect 3741 8120 3742 8440
rect 4062 8120 4063 8440
rect 3741 8119 4063 8120
rect 3318 7772 3422 8068
rect 2729 7720 3051 7721
rect 2729 7400 2730 7720
rect 3050 7400 3051 7720
rect 2729 7399 3051 7400
rect 2306 7052 2410 7348
rect 1717 7000 2039 7001
rect 1717 6680 1718 7000
rect 2038 6680 2039 7000
rect 1717 6679 2039 6680
rect 1294 6332 1398 6628
rect 705 6280 1027 6281
rect 705 5960 706 6280
rect 1026 5960 1027 6280
rect 705 5959 1027 5960
rect 282 5612 386 5908
rect -307 5560 15 5561
rect -307 5240 -306 5560
rect 14 5240 15 5560
rect -307 5239 15 5240
rect -730 4892 -626 5188
rect -1319 4840 -997 4841
rect -1319 4520 -1318 4840
rect -998 4520 -997 4840
rect -1319 4519 -997 4520
rect -1742 4172 -1638 4468
rect -2331 4120 -2009 4121
rect -2331 3800 -2330 4120
rect -2010 3800 -2009 4120
rect -2331 3799 -2009 3800
rect -2754 3452 -2650 3748
rect -3343 3400 -3021 3401
rect -3343 3080 -3342 3400
rect -3022 3080 -3021 3400
rect -3343 3079 -3021 3080
rect -3766 2732 -3662 3028
rect -4355 2680 -4033 2681
rect -4355 2360 -4354 2680
rect -4034 2360 -4033 2680
rect -4355 2359 -4033 2360
rect -4778 2012 -4674 2308
rect -5367 1960 -5045 1961
rect -5367 1640 -5366 1960
rect -5046 1640 -5045 1960
rect -5367 1639 -5045 1640
rect -5790 1292 -5686 1588
rect -6379 1240 -6057 1241
rect -6379 920 -6378 1240
rect -6058 920 -6057 1240
rect -6379 919 -6057 920
rect -6802 572 -6698 868
rect -7391 520 -7069 521
rect -7391 200 -7390 520
rect -7070 200 -7069 520
rect -7391 199 -7069 200
rect -7282 -199 -7178 199
rect -6802 148 -6782 572
rect -6718 148 -6698 572
rect -6270 521 -6166 919
rect -5790 868 -5770 1292
rect -5706 868 -5686 1292
rect -5258 1241 -5154 1639
rect -4778 1588 -4758 2012
rect -4694 1588 -4674 2012
rect -4246 1961 -4142 2359
rect -3766 2308 -3746 2732
rect -3682 2308 -3662 2732
rect -3234 2681 -3130 3079
rect -2754 3028 -2734 3452
rect -2670 3028 -2650 3452
rect -2222 3401 -2118 3799
rect -1742 3748 -1722 4172
rect -1658 3748 -1638 4172
rect -1210 4121 -1106 4519
rect -730 4468 -710 4892
rect -646 4468 -626 4892
rect -198 4841 -94 5239
rect 282 5188 302 5612
rect 366 5188 386 5612
rect 814 5561 918 5959
rect 1294 5908 1314 6332
rect 1378 5908 1398 6332
rect 1826 6281 1930 6679
rect 2306 6628 2326 7052
rect 2390 6628 2410 7052
rect 2838 7001 2942 7399
rect 3318 7348 3338 7772
rect 3402 7348 3422 7772
rect 3850 7721 3954 8119
rect 4330 8068 4350 8492
rect 4414 8068 4434 8492
rect 4862 8441 4966 8839
rect 5342 8788 5362 9212
rect 5426 8788 5446 9212
rect 5874 9161 5978 9559
rect 6354 9508 6374 9932
rect 6438 9508 6458 9932
rect 6886 9881 6990 10279
rect 7366 10228 7386 10652
rect 7450 10228 7470 10652
rect 7366 9932 7470 10228
rect 6777 9880 7099 9881
rect 6777 9560 6778 9880
rect 7098 9560 7099 9880
rect 6777 9559 7099 9560
rect 6354 9212 6458 9508
rect 5765 9160 6087 9161
rect 5765 8840 5766 9160
rect 6086 8840 6087 9160
rect 5765 8839 6087 8840
rect 5342 8492 5446 8788
rect 4753 8440 5075 8441
rect 4753 8120 4754 8440
rect 5074 8120 5075 8440
rect 4753 8119 5075 8120
rect 4330 7772 4434 8068
rect 3741 7720 4063 7721
rect 3741 7400 3742 7720
rect 4062 7400 4063 7720
rect 3741 7399 4063 7400
rect 3318 7052 3422 7348
rect 2729 7000 3051 7001
rect 2729 6680 2730 7000
rect 3050 6680 3051 7000
rect 2729 6679 3051 6680
rect 2306 6332 2410 6628
rect 1717 6280 2039 6281
rect 1717 5960 1718 6280
rect 2038 5960 2039 6280
rect 1717 5959 2039 5960
rect 1294 5612 1398 5908
rect 705 5560 1027 5561
rect 705 5240 706 5560
rect 1026 5240 1027 5560
rect 705 5239 1027 5240
rect 282 4892 386 5188
rect -307 4840 15 4841
rect -307 4520 -306 4840
rect 14 4520 15 4840
rect -307 4519 15 4520
rect -730 4172 -626 4468
rect -1319 4120 -997 4121
rect -1319 3800 -1318 4120
rect -998 3800 -997 4120
rect -1319 3799 -997 3800
rect -1742 3452 -1638 3748
rect -2331 3400 -2009 3401
rect -2331 3080 -2330 3400
rect -2010 3080 -2009 3400
rect -2331 3079 -2009 3080
rect -2754 2732 -2650 3028
rect -3343 2680 -3021 2681
rect -3343 2360 -3342 2680
rect -3022 2360 -3021 2680
rect -3343 2359 -3021 2360
rect -3766 2012 -3662 2308
rect -4355 1960 -4033 1961
rect -4355 1640 -4354 1960
rect -4034 1640 -4033 1960
rect -4355 1639 -4033 1640
rect -4778 1292 -4674 1588
rect -5367 1240 -5045 1241
rect -5367 920 -5366 1240
rect -5046 920 -5045 1240
rect -5367 919 -5045 920
rect -5790 572 -5686 868
rect -6379 520 -6057 521
rect -6379 200 -6378 520
rect -6058 200 -6057 520
rect -6379 199 -6057 200
rect -6802 -148 -6698 148
rect -7391 -200 -7069 -199
rect -7391 -520 -7390 -200
rect -7070 -520 -7069 -200
rect -7391 -521 -7069 -520
rect -7282 -919 -7178 -521
rect -6802 -572 -6782 -148
rect -6718 -572 -6698 -148
rect -6270 -199 -6166 199
rect -5790 148 -5770 572
rect -5706 148 -5686 572
rect -5258 521 -5154 919
rect -4778 868 -4758 1292
rect -4694 868 -4674 1292
rect -4246 1241 -4142 1639
rect -3766 1588 -3746 2012
rect -3682 1588 -3662 2012
rect -3234 1961 -3130 2359
rect -2754 2308 -2734 2732
rect -2670 2308 -2650 2732
rect -2222 2681 -2118 3079
rect -1742 3028 -1722 3452
rect -1658 3028 -1638 3452
rect -1210 3401 -1106 3799
rect -730 3748 -710 4172
rect -646 3748 -626 4172
rect -198 4121 -94 4519
rect 282 4468 302 4892
rect 366 4468 386 4892
rect 814 4841 918 5239
rect 1294 5188 1314 5612
rect 1378 5188 1398 5612
rect 1826 5561 1930 5959
rect 2306 5908 2326 6332
rect 2390 5908 2410 6332
rect 2838 6281 2942 6679
rect 3318 6628 3338 7052
rect 3402 6628 3422 7052
rect 3850 7001 3954 7399
rect 4330 7348 4350 7772
rect 4414 7348 4434 7772
rect 4862 7721 4966 8119
rect 5342 8068 5362 8492
rect 5426 8068 5446 8492
rect 5874 8441 5978 8839
rect 6354 8788 6374 9212
rect 6438 8788 6458 9212
rect 6886 9161 6990 9559
rect 7366 9508 7386 9932
rect 7450 9508 7470 9932
rect 7366 9212 7470 9508
rect 6777 9160 7099 9161
rect 6777 8840 6778 9160
rect 7098 8840 7099 9160
rect 6777 8839 7099 8840
rect 6354 8492 6458 8788
rect 5765 8440 6087 8441
rect 5765 8120 5766 8440
rect 6086 8120 6087 8440
rect 5765 8119 6087 8120
rect 5342 7772 5446 8068
rect 4753 7720 5075 7721
rect 4753 7400 4754 7720
rect 5074 7400 5075 7720
rect 4753 7399 5075 7400
rect 4330 7052 4434 7348
rect 3741 7000 4063 7001
rect 3741 6680 3742 7000
rect 4062 6680 4063 7000
rect 3741 6679 4063 6680
rect 3318 6332 3422 6628
rect 2729 6280 3051 6281
rect 2729 5960 2730 6280
rect 3050 5960 3051 6280
rect 2729 5959 3051 5960
rect 2306 5612 2410 5908
rect 1717 5560 2039 5561
rect 1717 5240 1718 5560
rect 2038 5240 2039 5560
rect 1717 5239 2039 5240
rect 1294 4892 1398 5188
rect 705 4840 1027 4841
rect 705 4520 706 4840
rect 1026 4520 1027 4840
rect 705 4519 1027 4520
rect 282 4172 386 4468
rect -307 4120 15 4121
rect -307 3800 -306 4120
rect 14 3800 15 4120
rect -307 3799 15 3800
rect -730 3452 -626 3748
rect -1319 3400 -997 3401
rect -1319 3080 -1318 3400
rect -998 3080 -997 3400
rect -1319 3079 -997 3080
rect -1742 2732 -1638 3028
rect -2331 2680 -2009 2681
rect -2331 2360 -2330 2680
rect -2010 2360 -2009 2680
rect -2331 2359 -2009 2360
rect -2754 2012 -2650 2308
rect -3343 1960 -3021 1961
rect -3343 1640 -3342 1960
rect -3022 1640 -3021 1960
rect -3343 1639 -3021 1640
rect -3766 1292 -3662 1588
rect -4355 1240 -4033 1241
rect -4355 920 -4354 1240
rect -4034 920 -4033 1240
rect -4355 919 -4033 920
rect -4778 572 -4674 868
rect -5367 520 -5045 521
rect -5367 200 -5366 520
rect -5046 200 -5045 520
rect -5367 199 -5045 200
rect -5790 -148 -5686 148
rect -6379 -200 -6057 -199
rect -6379 -520 -6378 -200
rect -6058 -520 -6057 -200
rect -6379 -521 -6057 -520
rect -6802 -868 -6698 -572
rect -7391 -920 -7069 -919
rect -7391 -1240 -7390 -920
rect -7070 -1240 -7069 -920
rect -7391 -1241 -7069 -1240
rect -7282 -1639 -7178 -1241
rect -6802 -1292 -6782 -868
rect -6718 -1292 -6698 -868
rect -6270 -919 -6166 -521
rect -5790 -572 -5770 -148
rect -5706 -572 -5686 -148
rect -5258 -199 -5154 199
rect -4778 148 -4758 572
rect -4694 148 -4674 572
rect -4246 521 -4142 919
rect -3766 868 -3746 1292
rect -3682 868 -3662 1292
rect -3234 1241 -3130 1639
rect -2754 1588 -2734 2012
rect -2670 1588 -2650 2012
rect -2222 1961 -2118 2359
rect -1742 2308 -1722 2732
rect -1658 2308 -1638 2732
rect -1210 2681 -1106 3079
rect -730 3028 -710 3452
rect -646 3028 -626 3452
rect -198 3401 -94 3799
rect 282 3748 302 4172
rect 366 3748 386 4172
rect 814 4121 918 4519
rect 1294 4468 1314 4892
rect 1378 4468 1398 4892
rect 1826 4841 1930 5239
rect 2306 5188 2326 5612
rect 2390 5188 2410 5612
rect 2838 5561 2942 5959
rect 3318 5908 3338 6332
rect 3402 5908 3422 6332
rect 3850 6281 3954 6679
rect 4330 6628 4350 7052
rect 4414 6628 4434 7052
rect 4862 7001 4966 7399
rect 5342 7348 5362 7772
rect 5426 7348 5446 7772
rect 5874 7721 5978 8119
rect 6354 8068 6374 8492
rect 6438 8068 6458 8492
rect 6886 8441 6990 8839
rect 7366 8788 7386 9212
rect 7450 8788 7470 9212
rect 7366 8492 7470 8788
rect 6777 8440 7099 8441
rect 6777 8120 6778 8440
rect 7098 8120 7099 8440
rect 6777 8119 7099 8120
rect 6354 7772 6458 8068
rect 5765 7720 6087 7721
rect 5765 7400 5766 7720
rect 6086 7400 6087 7720
rect 5765 7399 6087 7400
rect 5342 7052 5446 7348
rect 4753 7000 5075 7001
rect 4753 6680 4754 7000
rect 5074 6680 5075 7000
rect 4753 6679 5075 6680
rect 4330 6332 4434 6628
rect 3741 6280 4063 6281
rect 3741 5960 3742 6280
rect 4062 5960 4063 6280
rect 3741 5959 4063 5960
rect 3318 5612 3422 5908
rect 2729 5560 3051 5561
rect 2729 5240 2730 5560
rect 3050 5240 3051 5560
rect 2729 5239 3051 5240
rect 2306 4892 2410 5188
rect 1717 4840 2039 4841
rect 1717 4520 1718 4840
rect 2038 4520 2039 4840
rect 1717 4519 2039 4520
rect 1294 4172 1398 4468
rect 705 4120 1027 4121
rect 705 3800 706 4120
rect 1026 3800 1027 4120
rect 705 3799 1027 3800
rect 282 3452 386 3748
rect -307 3400 15 3401
rect -307 3080 -306 3400
rect 14 3080 15 3400
rect -307 3079 15 3080
rect -730 2732 -626 3028
rect -1319 2680 -997 2681
rect -1319 2360 -1318 2680
rect -998 2360 -997 2680
rect -1319 2359 -997 2360
rect -1742 2012 -1638 2308
rect -2331 1960 -2009 1961
rect -2331 1640 -2330 1960
rect -2010 1640 -2009 1960
rect -2331 1639 -2009 1640
rect -2754 1292 -2650 1588
rect -3343 1240 -3021 1241
rect -3343 920 -3342 1240
rect -3022 920 -3021 1240
rect -3343 919 -3021 920
rect -3766 572 -3662 868
rect -4355 520 -4033 521
rect -4355 200 -4354 520
rect -4034 200 -4033 520
rect -4355 199 -4033 200
rect -4778 -148 -4674 148
rect -5367 -200 -5045 -199
rect -5367 -520 -5366 -200
rect -5046 -520 -5045 -200
rect -5367 -521 -5045 -520
rect -5790 -868 -5686 -572
rect -6379 -920 -6057 -919
rect -6379 -1240 -6378 -920
rect -6058 -1240 -6057 -920
rect -6379 -1241 -6057 -1240
rect -6802 -1588 -6698 -1292
rect -7391 -1640 -7069 -1639
rect -7391 -1960 -7390 -1640
rect -7070 -1960 -7069 -1640
rect -7391 -1961 -7069 -1960
rect -7282 -2359 -7178 -1961
rect -6802 -2012 -6782 -1588
rect -6718 -2012 -6698 -1588
rect -6270 -1639 -6166 -1241
rect -5790 -1292 -5770 -868
rect -5706 -1292 -5686 -868
rect -5258 -919 -5154 -521
rect -4778 -572 -4758 -148
rect -4694 -572 -4674 -148
rect -4246 -199 -4142 199
rect -3766 148 -3746 572
rect -3682 148 -3662 572
rect -3234 521 -3130 919
rect -2754 868 -2734 1292
rect -2670 868 -2650 1292
rect -2222 1241 -2118 1639
rect -1742 1588 -1722 2012
rect -1658 1588 -1638 2012
rect -1210 1961 -1106 2359
rect -730 2308 -710 2732
rect -646 2308 -626 2732
rect -198 2681 -94 3079
rect 282 3028 302 3452
rect 366 3028 386 3452
rect 814 3401 918 3799
rect 1294 3748 1314 4172
rect 1378 3748 1398 4172
rect 1826 4121 1930 4519
rect 2306 4468 2326 4892
rect 2390 4468 2410 4892
rect 2838 4841 2942 5239
rect 3318 5188 3338 5612
rect 3402 5188 3422 5612
rect 3850 5561 3954 5959
rect 4330 5908 4350 6332
rect 4414 5908 4434 6332
rect 4862 6281 4966 6679
rect 5342 6628 5362 7052
rect 5426 6628 5446 7052
rect 5874 7001 5978 7399
rect 6354 7348 6374 7772
rect 6438 7348 6458 7772
rect 6886 7721 6990 8119
rect 7366 8068 7386 8492
rect 7450 8068 7470 8492
rect 7366 7772 7470 8068
rect 6777 7720 7099 7721
rect 6777 7400 6778 7720
rect 7098 7400 7099 7720
rect 6777 7399 7099 7400
rect 6354 7052 6458 7348
rect 5765 7000 6087 7001
rect 5765 6680 5766 7000
rect 6086 6680 6087 7000
rect 5765 6679 6087 6680
rect 5342 6332 5446 6628
rect 4753 6280 5075 6281
rect 4753 5960 4754 6280
rect 5074 5960 5075 6280
rect 4753 5959 5075 5960
rect 4330 5612 4434 5908
rect 3741 5560 4063 5561
rect 3741 5240 3742 5560
rect 4062 5240 4063 5560
rect 3741 5239 4063 5240
rect 3318 4892 3422 5188
rect 2729 4840 3051 4841
rect 2729 4520 2730 4840
rect 3050 4520 3051 4840
rect 2729 4519 3051 4520
rect 2306 4172 2410 4468
rect 1717 4120 2039 4121
rect 1717 3800 1718 4120
rect 2038 3800 2039 4120
rect 1717 3799 2039 3800
rect 1294 3452 1398 3748
rect 705 3400 1027 3401
rect 705 3080 706 3400
rect 1026 3080 1027 3400
rect 705 3079 1027 3080
rect 282 2732 386 3028
rect -307 2680 15 2681
rect -307 2360 -306 2680
rect 14 2360 15 2680
rect -307 2359 15 2360
rect -730 2012 -626 2308
rect -1319 1960 -997 1961
rect -1319 1640 -1318 1960
rect -998 1640 -997 1960
rect -1319 1639 -997 1640
rect -1742 1292 -1638 1588
rect -2331 1240 -2009 1241
rect -2331 920 -2330 1240
rect -2010 920 -2009 1240
rect -2331 919 -2009 920
rect -2754 572 -2650 868
rect -3343 520 -3021 521
rect -3343 200 -3342 520
rect -3022 200 -3021 520
rect -3343 199 -3021 200
rect -3766 -148 -3662 148
rect -4355 -200 -4033 -199
rect -4355 -520 -4354 -200
rect -4034 -520 -4033 -200
rect -4355 -521 -4033 -520
rect -4778 -868 -4674 -572
rect -5367 -920 -5045 -919
rect -5367 -1240 -5366 -920
rect -5046 -1240 -5045 -920
rect -5367 -1241 -5045 -1240
rect -5790 -1588 -5686 -1292
rect -6379 -1640 -6057 -1639
rect -6379 -1960 -6378 -1640
rect -6058 -1960 -6057 -1640
rect -6379 -1961 -6057 -1960
rect -6802 -2308 -6698 -2012
rect -7391 -2360 -7069 -2359
rect -7391 -2680 -7390 -2360
rect -7070 -2680 -7069 -2360
rect -7391 -2681 -7069 -2680
rect -7282 -3079 -7178 -2681
rect -6802 -2732 -6782 -2308
rect -6718 -2732 -6698 -2308
rect -6270 -2359 -6166 -1961
rect -5790 -2012 -5770 -1588
rect -5706 -2012 -5686 -1588
rect -5258 -1639 -5154 -1241
rect -4778 -1292 -4758 -868
rect -4694 -1292 -4674 -868
rect -4246 -919 -4142 -521
rect -3766 -572 -3746 -148
rect -3682 -572 -3662 -148
rect -3234 -199 -3130 199
rect -2754 148 -2734 572
rect -2670 148 -2650 572
rect -2222 521 -2118 919
rect -1742 868 -1722 1292
rect -1658 868 -1638 1292
rect -1210 1241 -1106 1639
rect -730 1588 -710 2012
rect -646 1588 -626 2012
rect -198 1961 -94 2359
rect 282 2308 302 2732
rect 366 2308 386 2732
rect 814 2681 918 3079
rect 1294 3028 1314 3452
rect 1378 3028 1398 3452
rect 1826 3401 1930 3799
rect 2306 3748 2326 4172
rect 2390 3748 2410 4172
rect 2838 4121 2942 4519
rect 3318 4468 3338 4892
rect 3402 4468 3422 4892
rect 3850 4841 3954 5239
rect 4330 5188 4350 5612
rect 4414 5188 4434 5612
rect 4862 5561 4966 5959
rect 5342 5908 5362 6332
rect 5426 5908 5446 6332
rect 5874 6281 5978 6679
rect 6354 6628 6374 7052
rect 6438 6628 6458 7052
rect 6886 7001 6990 7399
rect 7366 7348 7386 7772
rect 7450 7348 7470 7772
rect 7366 7052 7470 7348
rect 6777 7000 7099 7001
rect 6777 6680 6778 7000
rect 7098 6680 7099 7000
rect 6777 6679 7099 6680
rect 6354 6332 6458 6628
rect 5765 6280 6087 6281
rect 5765 5960 5766 6280
rect 6086 5960 6087 6280
rect 5765 5959 6087 5960
rect 5342 5612 5446 5908
rect 4753 5560 5075 5561
rect 4753 5240 4754 5560
rect 5074 5240 5075 5560
rect 4753 5239 5075 5240
rect 4330 4892 4434 5188
rect 3741 4840 4063 4841
rect 3741 4520 3742 4840
rect 4062 4520 4063 4840
rect 3741 4519 4063 4520
rect 3318 4172 3422 4468
rect 2729 4120 3051 4121
rect 2729 3800 2730 4120
rect 3050 3800 3051 4120
rect 2729 3799 3051 3800
rect 2306 3452 2410 3748
rect 1717 3400 2039 3401
rect 1717 3080 1718 3400
rect 2038 3080 2039 3400
rect 1717 3079 2039 3080
rect 1294 2732 1398 3028
rect 705 2680 1027 2681
rect 705 2360 706 2680
rect 1026 2360 1027 2680
rect 705 2359 1027 2360
rect 282 2012 386 2308
rect -307 1960 15 1961
rect -307 1640 -306 1960
rect 14 1640 15 1960
rect -307 1639 15 1640
rect -730 1292 -626 1588
rect -1319 1240 -997 1241
rect -1319 920 -1318 1240
rect -998 920 -997 1240
rect -1319 919 -997 920
rect -1742 572 -1638 868
rect -2331 520 -2009 521
rect -2331 200 -2330 520
rect -2010 200 -2009 520
rect -2331 199 -2009 200
rect -2754 -148 -2650 148
rect -3343 -200 -3021 -199
rect -3343 -520 -3342 -200
rect -3022 -520 -3021 -200
rect -3343 -521 -3021 -520
rect -3766 -868 -3662 -572
rect -4355 -920 -4033 -919
rect -4355 -1240 -4354 -920
rect -4034 -1240 -4033 -920
rect -4355 -1241 -4033 -1240
rect -4778 -1588 -4674 -1292
rect -5367 -1640 -5045 -1639
rect -5367 -1960 -5366 -1640
rect -5046 -1960 -5045 -1640
rect -5367 -1961 -5045 -1960
rect -5790 -2308 -5686 -2012
rect -6379 -2360 -6057 -2359
rect -6379 -2680 -6378 -2360
rect -6058 -2680 -6057 -2360
rect -6379 -2681 -6057 -2680
rect -6802 -3028 -6698 -2732
rect -7391 -3080 -7069 -3079
rect -7391 -3400 -7390 -3080
rect -7070 -3400 -7069 -3080
rect -7391 -3401 -7069 -3400
rect -7282 -3799 -7178 -3401
rect -6802 -3452 -6782 -3028
rect -6718 -3452 -6698 -3028
rect -6270 -3079 -6166 -2681
rect -5790 -2732 -5770 -2308
rect -5706 -2732 -5686 -2308
rect -5258 -2359 -5154 -1961
rect -4778 -2012 -4758 -1588
rect -4694 -2012 -4674 -1588
rect -4246 -1639 -4142 -1241
rect -3766 -1292 -3746 -868
rect -3682 -1292 -3662 -868
rect -3234 -919 -3130 -521
rect -2754 -572 -2734 -148
rect -2670 -572 -2650 -148
rect -2222 -199 -2118 199
rect -1742 148 -1722 572
rect -1658 148 -1638 572
rect -1210 521 -1106 919
rect -730 868 -710 1292
rect -646 868 -626 1292
rect -198 1241 -94 1639
rect 282 1588 302 2012
rect 366 1588 386 2012
rect 814 1961 918 2359
rect 1294 2308 1314 2732
rect 1378 2308 1398 2732
rect 1826 2681 1930 3079
rect 2306 3028 2326 3452
rect 2390 3028 2410 3452
rect 2838 3401 2942 3799
rect 3318 3748 3338 4172
rect 3402 3748 3422 4172
rect 3850 4121 3954 4519
rect 4330 4468 4350 4892
rect 4414 4468 4434 4892
rect 4862 4841 4966 5239
rect 5342 5188 5362 5612
rect 5426 5188 5446 5612
rect 5874 5561 5978 5959
rect 6354 5908 6374 6332
rect 6438 5908 6458 6332
rect 6886 6281 6990 6679
rect 7366 6628 7386 7052
rect 7450 6628 7470 7052
rect 7366 6332 7470 6628
rect 6777 6280 7099 6281
rect 6777 5960 6778 6280
rect 7098 5960 7099 6280
rect 6777 5959 7099 5960
rect 6354 5612 6458 5908
rect 5765 5560 6087 5561
rect 5765 5240 5766 5560
rect 6086 5240 6087 5560
rect 5765 5239 6087 5240
rect 5342 4892 5446 5188
rect 4753 4840 5075 4841
rect 4753 4520 4754 4840
rect 5074 4520 5075 4840
rect 4753 4519 5075 4520
rect 4330 4172 4434 4468
rect 3741 4120 4063 4121
rect 3741 3800 3742 4120
rect 4062 3800 4063 4120
rect 3741 3799 4063 3800
rect 3318 3452 3422 3748
rect 2729 3400 3051 3401
rect 2729 3080 2730 3400
rect 3050 3080 3051 3400
rect 2729 3079 3051 3080
rect 2306 2732 2410 3028
rect 1717 2680 2039 2681
rect 1717 2360 1718 2680
rect 2038 2360 2039 2680
rect 1717 2359 2039 2360
rect 1294 2012 1398 2308
rect 705 1960 1027 1961
rect 705 1640 706 1960
rect 1026 1640 1027 1960
rect 705 1639 1027 1640
rect 282 1292 386 1588
rect -307 1240 15 1241
rect -307 920 -306 1240
rect 14 920 15 1240
rect -307 919 15 920
rect -730 572 -626 868
rect -1319 520 -997 521
rect -1319 200 -1318 520
rect -998 200 -997 520
rect -1319 199 -997 200
rect -1742 -148 -1638 148
rect -2331 -200 -2009 -199
rect -2331 -520 -2330 -200
rect -2010 -520 -2009 -200
rect -2331 -521 -2009 -520
rect -2754 -868 -2650 -572
rect -3343 -920 -3021 -919
rect -3343 -1240 -3342 -920
rect -3022 -1240 -3021 -920
rect -3343 -1241 -3021 -1240
rect -3766 -1588 -3662 -1292
rect -4355 -1640 -4033 -1639
rect -4355 -1960 -4354 -1640
rect -4034 -1960 -4033 -1640
rect -4355 -1961 -4033 -1960
rect -4778 -2308 -4674 -2012
rect -5367 -2360 -5045 -2359
rect -5367 -2680 -5366 -2360
rect -5046 -2680 -5045 -2360
rect -5367 -2681 -5045 -2680
rect -5790 -3028 -5686 -2732
rect -6379 -3080 -6057 -3079
rect -6379 -3400 -6378 -3080
rect -6058 -3400 -6057 -3080
rect -6379 -3401 -6057 -3400
rect -6802 -3748 -6698 -3452
rect -7391 -3800 -7069 -3799
rect -7391 -4120 -7390 -3800
rect -7070 -4120 -7069 -3800
rect -7391 -4121 -7069 -4120
rect -7282 -4519 -7178 -4121
rect -6802 -4172 -6782 -3748
rect -6718 -4172 -6698 -3748
rect -6270 -3799 -6166 -3401
rect -5790 -3452 -5770 -3028
rect -5706 -3452 -5686 -3028
rect -5258 -3079 -5154 -2681
rect -4778 -2732 -4758 -2308
rect -4694 -2732 -4674 -2308
rect -4246 -2359 -4142 -1961
rect -3766 -2012 -3746 -1588
rect -3682 -2012 -3662 -1588
rect -3234 -1639 -3130 -1241
rect -2754 -1292 -2734 -868
rect -2670 -1292 -2650 -868
rect -2222 -919 -2118 -521
rect -1742 -572 -1722 -148
rect -1658 -572 -1638 -148
rect -1210 -199 -1106 199
rect -730 148 -710 572
rect -646 148 -626 572
rect -198 521 -94 919
rect 282 868 302 1292
rect 366 868 386 1292
rect 814 1241 918 1639
rect 1294 1588 1314 2012
rect 1378 1588 1398 2012
rect 1826 1961 1930 2359
rect 2306 2308 2326 2732
rect 2390 2308 2410 2732
rect 2838 2681 2942 3079
rect 3318 3028 3338 3452
rect 3402 3028 3422 3452
rect 3850 3401 3954 3799
rect 4330 3748 4350 4172
rect 4414 3748 4434 4172
rect 4862 4121 4966 4519
rect 5342 4468 5362 4892
rect 5426 4468 5446 4892
rect 5874 4841 5978 5239
rect 6354 5188 6374 5612
rect 6438 5188 6458 5612
rect 6886 5561 6990 5959
rect 7366 5908 7386 6332
rect 7450 5908 7470 6332
rect 7366 5612 7470 5908
rect 6777 5560 7099 5561
rect 6777 5240 6778 5560
rect 7098 5240 7099 5560
rect 6777 5239 7099 5240
rect 6354 4892 6458 5188
rect 5765 4840 6087 4841
rect 5765 4520 5766 4840
rect 6086 4520 6087 4840
rect 5765 4519 6087 4520
rect 5342 4172 5446 4468
rect 4753 4120 5075 4121
rect 4753 3800 4754 4120
rect 5074 3800 5075 4120
rect 4753 3799 5075 3800
rect 4330 3452 4434 3748
rect 3741 3400 4063 3401
rect 3741 3080 3742 3400
rect 4062 3080 4063 3400
rect 3741 3079 4063 3080
rect 3318 2732 3422 3028
rect 2729 2680 3051 2681
rect 2729 2360 2730 2680
rect 3050 2360 3051 2680
rect 2729 2359 3051 2360
rect 2306 2012 2410 2308
rect 1717 1960 2039 1961
rect 1717 1640 1718 1960
rect 2038 1640 2039 1960
rect 1717 1639 2039 1640
rect 1294 1292 1398 1588
rect 705 1240 1027 1241
rect 705 920 706 1240
rect 1026 920 1027 1240
rect 705 919 1027 920
rect 282 572 386 868
rect -307 520 15 521
rect -307 200 -306 520
rect 14 200 15 520
rect -307 199 15 200
rect -730 -148 -626 148
rect -1319 -200 -997 -199
rect -1319 -520 -1318 -200
rect -998 -520 -997 -200
rect -1319 -521 -997 -520
rect -1742 -868 -1638 -572
rect -2331 -920 -2009 -919
rect -2331 -1240 -2330 -920
rect -2010 -1240 -2009 -920
rect -2331 -1241 -2009 -1240
rect -2754 -1588 -2650 -1292
rect -3343 -1640 -3021 -1639
rect -3343 -1960 -3342 -1640
rect -3022 -1960 -3021 -1640
rect -3343 -1961 -3021 -1960
rect -3766 -2308 -3662 -2012
rect -4355 -2360 -4033 -2359
rect -4355 -2680 -4354 -2360
rect -4034 -2680 -4033 -2360
rect -4355 -2681 -4033 -2680
rect -4778 -3028 -4674 -2732
rect -5367 -3080 -5045 -3079
rect -5367 -3400 -5366 -3080
rect -5046 -3400 -5045 -3080
rect -5367 -3401 -5045 -3400
rect -5790 -3748 -5686 -3452
rect -6379 -3800 -6057 -3799
rect -6379 -4120 -6378 -3800
rect -6058 -4120 -6057 -3800
rect -6379 -4121 -6057 -4120
rect -6802 -4468 -6698 -4172
rect -7391 -4520 -7069 -4519
rect -7391 -4840 -7390 -4520
rect -7070 -4840 -7069 -4520
rect -7391 -4841 -7069 -4840
rect -7282 -5239 -7178 -4841
rect -6802 -4892 -6782 -4468
rect -6718 -4892 -6698 -4468
rect -6270 -4519 -6166 -4121
rect -5790 -4172 -5770 -3748
rect -5706 -4172 -5686 -3748
rect -5258 -3799 -5154 -3401
rect -4778 -3452 -4758 -3028
rect -4694 -3452 -4674 -3028
rect -4246 -3079 -4142 -2681
rect -3766 -2732 -3746 -2308
rect -3682 -2732 -3662 -2308
rect -3234 -2359 -3130 -1961
rect -2754 -2012 -2734 -1588
rect -2670 -2012 -2650 -1588
rect -2222 -1639 -2118 -1241
rect -1742 -1292 -1722 -868
rect -1658 -1292 -1638 -868
rect -1210 -919 -1106 -521
rect -730 -572 -710 -148
rect -646 -572 -626 -148
rect -198 -199 -94 199
rect 282 148 302 572
rect 366 148 386 572
rect 814 521 918 919
rect 1294 868 1314 1292
rect 1378 868 1398 1292
rect 1826 1241 1930 1639
rect 2306 1588 2326 2012
rect 2390 1588 2410 2012
rect 2838 1961 2942 2359
rect 3318 2308 3338 2732
rect 3402 2308 3422 2732
rect 3850 2681 3954 3079
rect 4330 3028 4350 3452
rect 4414 3028 4434 3452
rect 4862 3401 4966 3799
rect 5342 3748 5362 4172
rect 5426 3748 5446 4172
rect 5874 4121 5978 4519
rect 6354 4468 6374 4892
rect 6438 4468 6458 4892
rect 6886 4841 6990 5239
rect 7366 5188 7386 5612
rect 7450 5188 7470 5612
rect 7366 4892 7470 5188
rect 6777 4840 7099 4841
rect 6777 4520 6778 4840
rect 7098 4520 7099 4840
rect 6777 4519 7099 4520
rect 6354 4172 6458 4468
rect 5765 4120 6087 4121
rect 5765 3800 5766 4120
rect 6086 3800 6087 4120
rect 5765 3799 6087 3800
rect 5342 3452 5446 3748
rect 4753 3400 5075 3401
rect 4753 3080 4754 3400
rect 5074 3080 5075 3400
rect 4753 3079 5075 3080
rect 4330 2732 4434 3028
rect 3741 2680 4063 2681
rect 3741 2360 3742 2680
rect 4062 2360 4063 2680
rect 3741 2359 4063 2360
rect 3318 2012 3422 2308
rect 2729 1960 3051 1961
rect 2729 1640 2730 1960
rect 3050 1640 3051 1960
rect 2729 1639 3051 1640
rect 2306 1292 2410 1588
rect 1717 1240 2039 1241
rect 1717 920 1718 1240
rect 2038 920 2039 1240
rect 1717 919 2039 920
rect 1294 572 1398 868
rect 705 520 1027 521
rect 705 200 706 520
rect 1026 200 1027 520
rect 705 199 1027 200
rect 282 -148 386 148
rect -307 -200 15 -199
rect -307 -520 -306 -200
rect 14 -520 15 -200
rect -307 -521 15 -520
rect -730 -868 -626 -572
rect -1319 -920 -997 -919
rect -1319 -1240 -1318 -920
rect -998 -1240 -997 -920
rect -1319 -1241 -997 -1240
rect -1742 -1588 -1638 -1292
rect -2331 -1640 -2009 -1639
rect -2331 -1960 -2330 -1640
rect -2010 -1960 -2009 -1640
rect -2331 -1961 -2009 -1960
rect -2754 -2308 -2650 -2012
rect -3343 -2360 -3021 -2359
rect -3343 -2680 -3342 -2360
rect -3022 -2680 -3021 -2360
rect -3343 -2681 -3021 -2680
rect -3766 -3028 -3662 -2732
rect -4355 -3080 -4033 -3079
rect -4355 -3400 -4354 -3080
rect -4034 -3400 -4033 -3080
rect -4355 -3401 -4033 -3400
rect -4778 -3748 -4674 -3452
rect -5367 -3800 -5045 -3799
rect -5367 -4120 -5366 -3800
rect -5046 -4120 -5045 -3800
rect -5367 -4121 -5045 -4120
rect -5790 -4468 -5686 -4172
rect -6379 -4520 -6057 -4519
rect -6379 -4840 -6378 -4520
rect -6058 -4840 -6057 -4520
rect -6379 -4841 -6057 -4840
rect -6802 -5188 -6698 -4892
rect -7391 -5240 -7069 -5239
rect -7391 -5560 -7390 -5240
rect -7070 -5560 -7069 -5240
rect -7391 -5561 -7069 -5560
rect -7282 -5959 -7178 -5561
rect -6802 -5612 -6782 -5188
rect -6718 -5612 -6698 -5188
rect -6270 -5239 -6166 -4841
rect -5790 -4892 -5770 -4468
rect -5706 -4892 -5686 -4468
rect -5258 -4519 -5154 -4121
rect -4778 -4172 -4758 -3748
rect -4694 -4172 -4674 -3748
rect -4246 -3799 -4142 -3401
rect -3766 -3452 -3746 -3028
rect -3682 -3452 -3662 -3028
rect -3234 -3079 -3130 -2681
rect -2754 -2732 -2734 -2308
rect -2670 -2732 -2650 -2308
rect -2222 -2359 -2118 -1961
rect -1742 -2012 -1722 -1588
rect -1658 -2012 -1638 -1588
rect -1210 -1639 -1106 -1241
rect -730 -1292 -710 -868
rect -646 -1292 -626 -868
rect -198 -919 -94 -521
rect 282 -572 302 -148
rect 366 -572 386 -148
rect 814 -199 918 199
rect 1294 148 1314 572
rect 1378 148 1398 572
rect 1826 521 1930 919
rect 2306 868 2326 1292
rect 2390 868 2410 1292
rect 2838 1241 2942 1639
rect 3318 1588 3338 2012
rect 3402 1588 3422 2012
rect 3850 1961 3954 2359
rect 4330 2308 4350 2732
rect 4414 2308 4434 2732
rect 4862 2681 4966 3079
rect 5342 3028 5362 3452
rect 5426 3028 5446 3452
rect 5874 3401 5978 3799
rect 6354 3748 6374 4172
rect 6438 3748 6458 4172
rect 6886 4121 6990 4519
rect 7366 4468 7386 4892
rect 7450 4468 7470 4892
rect 7366 4172 7470 4468
rect 6777 4120 7099 4121
rect 6777 3800 6778 4120
rect 7098 3800 7099 4120
rect 6777 3799 7099 3800
rect 6354 3452 6458 3748
rect 5765 3400 6087 3401
rect 5765 3080 5766 3400
rect 6086 3080 6087 3400
rect 5765 3079 6087 3080
rect 5342 2732 5446 3028
rect 4753 2680 5075 2681
rect 4753 2360 4754 2680
rect 5074 2360 5075 2680
rect 4753 2359 5075 2360
rect 4330 2012 4434 2308
rect 3741 1960 4063 1961
rect 3741 1640 3742 1960
rect 4062 1640 4063 1960
rect 3741 1639 4063 1640
rect 3318 1292 3422 1588
rect 2729 1240 3051 1241
rect 2729 920 2730 1240
rect 3050 920 3051 1240
rect 2729 919 3051 920
rect 2306 572 2410 868
rect 1717 520 2039 521
rect 1717 200 1718 520
rect 2038 200 2039 520
rect 1717 199 2039 200
rect 1294 -148 1398 148
rect 705 -200 1027 -199
rect 705 -520 706 -200
rect 1026 -520 1027 -200
rect 705 -521 1027 -520
rect 282 -868 386 -572
rect -307 -920 15 -919
rect -307 -1240 -306 -920
rect 14 -1240 15 -920
rect -307 -1241 15 -1240
rect -730 -1588 -626 -1292
rect -1319 -1640 -997 -1639
rect -1319 -1960 -1318 -1640
rect -998 -1960 -997 -1640
rect -1319 -1961 -997 -1960
rect -1742 -2308 -1638 -2012
rect -2331 -2360 -2009 -2359
rect -2331 -2680 -2330 -2360
rect -2010 -2680 -2009 -2360
rect -2331 -2681 -2009 -2680
rect -2754 -3028 -2650 -2732
rect -3343 -3080 -3021 -3079
rect -3343 -3400 -3342 -3080
rect -3022 -3400 -3021 -3080
rect -3343 -3401 -3021 -3400
rect -3766 -3748 -3662 -3452
rect -4355 -3800 -4033 -3799
rect -4355 -4120 -4354 -3800
rect -4034 -4120 -4033 -3800
rect -4355 -4121 -4033 -4120
rect -4778 -4468 -4674 -4172
rect -5367 -4520 -5045 -4519
rect -5367 -4840 -5366 -4520
rect -5046 -4840 -5045 -4520
rect -5367 -4841 -5045 -4840
rect -5790 -5188 -5686 -4892
rect -6379 -5240 -6057 -5239
rect -6379 -5560 -6378 -5240
rect -6058 -5560 -6057 -5240
rect -6379 -5561 -6057 -5560
rect -6802 -5908 -6698 -5612
rect -7391 -5960 -7069 -5959
rect -7391 -6280 -7390 -5960
rect -7070 -6280 -7069 -5960
rect -7391 -6281 -7069 -6280
rect -7282 -6679 -7178 -6281
rect -6802 -6332 -6782 -5908
rect -6718 -6332 -6698 -5908
rect -6270 -5959 -6166 -5561
rect -5790 -5612 -5770 -5188
rect -5706 -5612 -5686 -5188
rect -5258 -5239 -5154 -4841
rect -4778 -4892 -4758 -4468
rect -4694 -4892 -4674 -4468
rect -4246 -4519 -4142 -4121
rect -3766 -4172 -3746 -3748
rect -3682 -4172 -3662 -3748
rect -3234 -3799 -3130 -3401
rect -2754 -3452 -2734 -3028
rect -2670 -3452 -2650 -3028
rect -2222 -3079 -2118 -2681
rect -1742 -2732 -1722 -2308
rect -1658 -2732 -1638 -2308
rect -1210 -2359 -1106 -1961
rect -730 -2012 -710 -1588
rect -646 -2012 -626 -1588
rect -198 -1639 -94 -1241
rect 282 -1292 302 -868
rect 366 -1292 386 -868
rect 814 -919 918 -521
rect 1294 -572 1314 -148
rect 1378 -572 1398 -148
rect 1826 -199 1930 199
rect 2306 148 2326 572
rect 2390 148 2410 572
rect 2838 521 2942 919
rect 3318 868 3338 1292
rect 3402 868 3422 1292
rect 3850 1241 3954 1639
rect 4330 1588 4350 2012
rect 4414 1588 4434 2012
rect 4862 1961 4966 2359
rect 5342 2308 5362 2732
rect 5426 2308 5446 2732
rect 5874 2681 5978 3079
rect 6354 3028 6374 3452
rect 6438 3028 6458 3452
rect 6886 3401 6990 3799
rect 7366 3748 7386 4172
rect 7450 3748 7470 4172
rect 7366 3452 7470 3748
rect 6777 3400 7099 3401
rect 6777 3080 6778 3400
rect 7098 3080 7099 3400
rect 6777 3079 7099 3080
rect 6354 2732 6458 3028
rect 5765 2680 6087 2681
rect 5765 2360 5766 2680
rect 6086 2360 6087 2680
rect 5765 2359 6087 2360
rect 5342 2012 5446 2308
rect 4753 1960 5075 1961
rect 4753 1640 4754 1960
rect 5074 1640 5075 1960
rect 4753 1639 5075 1640
rect 4330 1292 4434 1588
rect 3741 1240 4063 1241
rect 3741 920 3742 1240
rect 4062 920 4063 1240
rect 3741 919 4063 920
rect 3318 572 3422 868
rect 2729 520 3051 521
rect 2729 200 2730 520
rect 3050 200 3051 520
rect 2729 199 3051 200
rect 2306 -148 2410 148
rect 1717 -200 2039 -199
rect 1717 -520 1718 -200
rect 2038 -520 2039 -200
rect 1717 -521 2039 -520
rect 1294 -868 1398 -572
rect 705 -920 1027 -919
rect 705 -1240 706 -920
rect 1026 -1240 1027 -920
rect 705 -1241 1027 -1240
rect 282 -1588 386 -1292
rect -307 -1640 15 -1639
rect -307 -1960 -306 -1640
rect 14 -1960 15 -1640
rect -307 -1961 15 -1960
rect -730 -2308 -626 -2012
rect -1319 -2360 -997 -2359
rect -1319 -2680 -1318 -2360
rect -998 -2680 -997 -2360
rect -1319 -2681 -997 -2680
rect -1742 -3028 -1638 -2732
rect -2331 -3080 -2009 -3079
rect -2331 -3400 -2330 -3080
rect -2010 -3400 -2009 -3080
rect -2331 -3401 -2009 -3400
rect -2754 -3748 -2650 -3452
rect -3343 -3800 -3021 -3799
rect -3343 -4120 -3342 -3800
rect -3022 -4120 -3021 -3800
rect -3343 -4121 -3021 -4120
rect -3766 -4468 -3662 -4172
rect -4355 -4520 -4033 -4519
rect -4355 -4840 -4354 -4520
rect -4034 -4840 -4033 -4520
rect -4355 -4841 -4033 -4840
rect -4778 -5188 -4674 -4892
rect -5367 -5240 -5045 -5239
rect -5367 -5560 -5366 -5240
rect -5046 -5560 -5045 -5240
rect -5367 -5561 -5045 -5560
rect -5790 -5908 -5686 -5612
rect -6379 -5960 -6057 -5959
rect -6379 -6280 -6378 -5960
rect -6058 -6280 -6057 -5960
rect -6379 -6281 -6057 -6280
rect -6802 -6628 -6698 -6332
rect -7391 -6680 -7069 -6679
rect -7391 -7000 -7390 -6680
rect -7070 -7000 -7069 -6680
rect -7391 -7001 -7069 -7000
rect -7282 -7399 -7178 -7001
rect -6802 -7052 -6782 -6628
rect -6718 -7052 -6698 -6628
rect -6270 -6679 -6166 -6281
rect -5790 -6332 -5770 -5908
rect -5706 -6332 -5686 -5908
rect -5258 -5959 -5154 -5561
rect -4778 -5612 -4758 -5188
rect -4694 -5612 -4674 -5188
rect -4246 -5239 -4142 -4841
rect -3766 -4892 -3746 -4468
rect -3682 -4892 -3662 -4468
rect -3234 -4519 -3130 -4121
rect -2754 -4172 -2734 -3748
rect -2670 -4172 -2650 -3748
rect -2222 -3799 -2118 -3401
rect -1742 -3452 -1722 -3028
rect -1658 -3452 -1638 -3028
rect -1210 -3079 -1106 -2681
rect -730 -2732 -710 -2308
rect -646 -2732 -626 -2308
rect -198 -2359 -94 -1961
rect 282 -2012 302 -1588
rect 366 -2012 386 -1588
rect 814 -1639 918 -1241
rect 1294 -1292 1314 -868
rect 1378 -1292 1398 -868
rect 1826 -919 1930 -521
rect 2306 -572 2326 -148
rect 2390 -572 2410 -148
rect 2838 -199 2942 199
rect 3318 148 3338 572
rect 3402 148 3422 572
rect 3850 521 3954 919
rect 4330 868 4350 1292
rect 4414 868 4434 1292
rect 4862 1241 4966 1639
rect 5342 1588 5362 2012
rect 5426 1588 5446 2012
rect 5874 1961 5978 2359
rect 6354 2308 6374 2732
rect 6438 2308 6458 2732
rect 6886 2681 6990 3079
rect 7366 3028 7386 3452
rect 7450 3028 7470 3452
rect 7366 2732 7470 3028
rect 6777 2680 7099 2681
rect 6777 2360 6778 2680
rect 7098 2360 7099 2680
rect 6777 2359 7099 2360
rect 6354 2012 6458 2308
rect 5765 1960 6087 1961
rect 5765 1640 5766 1960
rect 6086 1640 6087 1960
rect 5765 1639 6087 1640
rect 5342 1292 5446 1588
rect 4753 1240 5075 1241
rect 4753 920 4754 1240
rect 5074 920 5075 1240
rect 4753 919 5075 920
rect 4330 572 4434 868
rect 3741 520 4063 521
rect 3741 200 3742 520
rect 4062 200 4063 520
rect 3741 199 4063 200
rect 3318 -148 3422 148
rect 2729 -200 3051 -199
rect 2729 -520 2730 -200
rect 3050 -520 3051 -200
rect 2729 -521 3051 -520
rect 2306 -868 2410 -572
rect 1717 -920 2039 -919
rect 1717 -1240 1718 -920
rect 2038 -1240 2039 -920
rect 1717 -1241 2039 -1240
rect 1294 -1588 1398 -1292
rect 705 -1640 1027 -1639
rect 705 -1960 706 -1640
rect 1026 -1960 1027 -1640
rect 705 -1961 1027 -1960
rect 282 -2308 386 -2012
rect -307 -2360 15 -2359
rect -307 -2680 -306 -2360
rect 14 -2680 15 -2360
rect -307 -2681 15 -2680
rect -730 -3028 -626 -2732
rect -1319 -3080 -997 -3079
rect -1319 -3400 -1318 -3080
rect -998 -3400 -997 -3080
rect -1319 -3401 -997 -3400
rect -1742 -3748 -1638 -3452
rect -2331 -3800 -2009 -3799
rect -2331 -4120 -2330 -3800
rect -2010 -4120 -2009 -3800
rect -2331 -4121 -2009 -4120
rect -2754 -4468 -2650 -4172
rect -3343 -4520 -3021 -4519
rect -3343 -4840 -3342 -4520
rect -3022 -4840 -3021 -4520
rect -3343 -4841 -3021 -4840
rect -3766 -5188 -3662 -4892
rect -4355 -5240 -4033 -5239
rect -4355 -5560 -4354 -5240
rect -4034 -5560 -4033 -5240
rect -4355 -5561 -4033 -5560
rect -4778 -5908 -4674 -5612
rect -5367 -5960 -5045 -5959
rect -5367 -6280 -5366 -5960
rect -5046 -6280 -5045 -5960
rect -5367 -6281 -5045 -6280
rect -5790 -6628 -5686 -6332
rect -6379 -6680 -6057 -6679
rect -6379 -7000 -6378 -6680
rect -6058 -7000 -6057 -6680
rect -6379 -7001 -6057 -7000
rect -6802 -7348 -6698 -7052
rect -7391 -7400 -7069 -7399
rect -7391 -7720 -7390 -7400
rect -7070 -7720 -7069 -7400
rect -7391 -7721 -7069 -7720
rect -7282 -8119 -7178 -7721
rect -6802 -7772 -6782 -7348
rect -6718 -7772 -6698 -7348
rect -6270 -7399 -6166 -7001
rect -5790 -7052 -5770 -6628
rect -5706 -7052 -5686 -6628
rect -5258 -6679 -5154 -6281
rect -4778 -6332 -4758 -5908
rect -4694 -6332 -4674 -5908
rect -4246 -5959 -4142 -5561
rect -3766 -5612 -3746 -5188
rect -3682 -5612 -3662 -5188
rect -3234 -5239 -3130 -4841
rect -2754 -4892 -2734 -4468
rect -2670 -4892 -2650 -4468
rect -2222 -4519 -2118 -4121
rect -1742 -4172 -1722 -3748
rect -1658 -4172 -1638 -3748
rect -1210 -3799 -1106 -3401
rect -730 -3452 -710 -3028
rect -646 -3452 -626 -3028
rect -198 -3079 -94 -2681
rect 282 -2732 302 -2308
rect 366 -2732 386 -2308
rect 814 -2359 918 -1961
rect 1294 -2012 1314 -1588
rect 1378 -2012 1398 -1588
rect 1826 -1639 1930 -1241
rect 2306 -1292 2326 -868
rect 2390 -1292 2410 -868
rect 2838 -919 2942 -521
rect 3318 -572 3338 -148
rect 3402 -572 3422 -148
rect 3850 -199 3954 199
rect 4330 148 4350 572
rect 4414 148 4434 572
rect 4862 521 4966 919
rect 5342 868 5362 1292
rect 5426 868 5446 1292
rect 5874 1241 5978 1639
rect 6354 1588 6374 2012
rect 6438 1588 6458 2012
rect 6886 1961 6990 2359
rect 7366 2308 7386 2732
rect 7450 2308 7470 2732
rect 7366 2012 7470 2308
rect 6777 1960 7099 1961
rect 6777 1640 6778 1960
rect 7098 1640 7099 1960
rect 6777 1639 7099 1640
rect 6354 1292 6458 1588
rect 5765 1240 6087 1241
rect 5765 920 5766 1240
rect 6086 920 6087 1240
rect 5765 919 6087 920
rect 5342 572 5446 868
rect 4753 520 5075 521
rect 4753 200 4754 520
rect 5074 200 5075 520
rect 4753 199 5075 200
rect 4330 -148 4434 148
rect 3741 -200 4063 -199
rect 3741 -520 3742 -200
rect 4062 -520 4063 -200
rect 3741 -521 4063 -520
rect 3318 -868 3422 -572
rect 2729 -920 3051 -919
rect 2729 -1240 2730 -920
rect 3050 -1240 3051 -920
rect 2729 -1241 3051 -1240
rect 2306 -1588 2410 -1292
rect 1717 -1640 2039 -1639
rect 1717 -1960 1718 -1640
rect 2038 -1960 2039 -1640
rect 1717 -1961 2039 -1960
rect 1294 -2308 1398 -2012
rect 705 -2360 1027 -2359
rect 705 -2680 706 -2360
rect 1026 -2680 1027 -2360
rect 705 -2681 1027 -2680
rect 282 -3028 386 -2732
rect -307 -3080 15 -3079
rect -307 -3400 -306 -3080
rect 14 -3400 15 -3080
rect -307 -3401 15 -3400
rect -730 -3748 -626 -3452
rect -1319 -3800 -997 -3799
rect -1319 -4120 -1318 -3800
rect -998 -4120 -997 -3800
rect -1319 -4121 -997 -4120
rect -1742 -4468 -1638 -4172
rect -2331 -4520 -2009 -4519
rect -2331 -4840 -2330 -4520
rect -2010 -4840 -2009 -4520
rect -2331 -4841 -2009 -4840
rect -2754 -5188 -2650 -4892
rect -3343 -5240 -3021 -5239
rect -3343 -5560 -3342 -5240
rect -3022 -5560 -3021 -5240
rect -3343 -5561 -3021 -5560
rect -3766 -5908 -3662 -5612
rect -4355 -5960 -4033 -5959
rect -4355 -6280 -4354 -5960
rect -4034 -6280 -4033 -5960
rect -4355 -6281 -4033 -6280
rect -4778 -6628 -4674 -6332
rect -5367 -6680 -5045 -6679
rect -5367 -7000 -5366 -6680
rect -5046 -7000 -5045 -6680
rect -5367 -7001 -5045 -7000
rect -5790 -7348 -5686 -7052
rect -6379 -7400 -6057 -7399
rect -6379 -7720 -6378 -7400
rect -6058 -7720 -6057 -7400
rect -6379 -7721 -6057 -7720
rect -6802 -8068 -6698 -7772
rect -7391 -8120 -7069 -8119
rect -7391 -8440 -7390 -8120
rect -7070 -8440 -7069 -8120
rect -7391 -8441 -7069 -8440
rect -7282 -8839 -7178 -8441
rect -6802 -8492 -6782 -8068
rect -6718 -8492 -6698 -8068
rect -6270 -8119 -6166 -7721
rect -5790 -7772 -5770 -7348
rect -5706 -7772 -5686 -7348
rect -5258 -7399 -5154 -7001
rect -4778 -7052 -4758 -6628
rect -4694 -7052 -4674 -6628
rect -4246 -6679 -4142 -6281
rect -3766 -6332 -3746 -5908
rect -3682 -6332 -3662 -5908
rect -3234 -5959 -3130 -5561
rect -2754 -5612 -2734 -5188
rect -2670 -5612 -2650 -5188
rect -2222 -5239 -2118 -4841
rect -1742 -4892 -1722 -4468
rect -1658 -4892 -1638 -4468
rect -1210 -4519 -1106 -4121
rect -730 -4172 -710 -3748
rect -646 -4172 -626 -3748
rect -198 -3799 -94 -3401
rect 282 -3452 302 -3028
rect 366 -3452 386 -3028
rect 814 -3079 918 -2681
rect 1294 -2732 1314 -2308
rect 1378 -2732 1398 -2308
rect 1826 -2359 1930 -1961
rect 2306 -2012 2326 -1588
rect 2390 -2012 2410 -1588
rect 2838 -1639 2942 -1241
rect 3318 -1292 3338 -868
rect 3402 -1292 3422 -868
rect 3850 -919 3954 -521
rect 4330 -572 4350 -148
rect 4414 -572 4434 -148
rect 4862 -199 4966 199
rect 5342 148 5362 572
rect 5426 148 5446 572
rect 5874 521 5978 919
rect 6354 868 6374 1292
rect 6438 868 6458 1292
rect 6886 1241 6990 1639
rect 7366 1588 7386 2012
rect 7450 1588 7470 2012
rect 7366 1292 7470 1588
rect 6777 1240 7099 1241
rect 6777 920 6778 1240
rect 7098 920 7099 1240
rect 6777 919 7099 920
rect 6354 572 6458 868
rect 5765 520 6087 521
rect 5765 200 5766 520
rect 6086 200 6087 520
rect 5765 199 6087 200
rect 5342 -148 5446 148
rect 4753 -200 5075 -199
rect 4753 -520 4754 -200
rect 5074 -520 5075 -200
rect 4753 -521 5075 -520
rect 4330 -868 4434 -572
rect 3741 -920 4063 -919
rect 3741 -1240 3742 -920
rect 4062 -1240 4063 -920
rect 3741 -1241 4063 -1240
rect 3318 -1588 3422 -1292
rect 2729 -1640 3051 -1639
rect 2729 -1960 2730 -1640
rect 3050 -1960 3051 -1640
rect 2729 -1961 3051 -1960
rect 2306 -2308 2410 -2012
rect 1717 -2360 2039 -2359
rect 1717 -2680 1718 -2360
rect 2038 -2680 2039 -2360
rect 1717 -2681 2039 -2680
rect 1294 -3028 1398 -2732
rect 705 -3080 1027 -3079
rect 705 -3400 706 -3080
rect 1026 -3400 1027 -3080
rect 705 -3401 1027 -3400
rect 282 -3748 386 -3452
rect -307 -3800 15 -3799
rect -307 -4120 -306 -3800
rect 14 -4120 15 -3800
rect -307 -4121 15 -4120
rect -730 -4468 -626 -4172
rect -1319 -4520 -997 -4519
rect -1319 -4840 -1318 -4520
rect -998 -4840 -997 -4520
rect -1319 -4841 -997 -4840
rect -1742 -5188 -1638 -4892
rect -2331 -5240 -2009 -5239
rect -2331 -5560 -2330 -5240
rect -2010 -5560 -2009 -5240
rect -2331 -5561 -2009 -5560
rect -2754 -5908 -2650 -5612
rect -3343 -5960 -3021 -5959
rect -3343 -6280 -3342 -5960
rect -3022 -6280 -3021 -5960
rect -3343 -6281 -3021 -6280
rect -3766 -6628 -3662 -6332
rect -4355 -6680 -4033 -6679
rect -4355 -7000 -4354 -6680
rect -4034 -7000 -4033 -6680
rect -4355 -7001 -4033 -7000
rect -4778 -7348 -4674 -7052
rect -5367 -7400 -5045 -7399
rect -5367 -7720 -5366 -7400
rect -5046 -7720 -5045 -7400
rect -5367 -7721 -5045 -7720
rect -5790 -8068 -5686 -7772
rect -6379 -8120 -6057 -8119
rect -6379 -8440 -6378 -8120
rect -6058 -8440 -6057 -8120
rect -6379 -8441 -6057 -8440
rect -6802 -8788 -6698 -8492
rect -7391 -8840 -7069 -8839
rect -7391 -9160 -7390 -8840
rect -7070 -9160 -7069 -8840
rect -7391 -9161 -7069 -9160
rect -7282 -9559 -7178 -9161
rect -6802 -9212 -6782 -8788
rect -6718 -9212 -6698 -8788
rect -6270 -8839 -6166 -8441
rect -5790 -8492 -5770 -8068
rect -5706 -8492 -5686 -8068
rect -5258 -8119 -5154 -7721
rect -4778 -7772 -4758 -7348
rect -4694 -7772 -4674 -7348
rect -4246 -7399 -4142 -7001
rect -3766 -7052 -3746 -6628
rect -3682 -7052 -3662 -6628
rect -3234 -6679 -3130 -6281
rect -2754 -6332 -2734 -5908
rect -2670 -6332 -2650 -5908
rect -2222 -5959 -2118 -5561
rect -1742 -5612 -1722 -5188
rect -1658 -5612 -1638 -5188
rect -1210 -5239 -1106 -4841
rect -730 -4892 -710 -4468
rect -646 -4892 -626 -4468
rect -198 -4519 -94 -4121
rect 282 -4172 302 -3748
rect 366 -4172 386 -3748
rect 814 -3799 918 -3401
rect 1294 -3452 1314 -3028
rect 1378 -3452 1398 -3028
rect 1826 -3079 1930 -2681
rect 2306 -2732 2326 -2308
rect 2390 -2732 2410 -2308
rect 2838 -2359 2942 -1961
rect 3318 -2012 3338 -1588
rect 3402 -2012 3422 -1588
rect 3850 -1639 3954 -1241
rect 4330 -1292 4350 -868
rect 4414 -1292 4434 -868
rect 4862 -919 4966 -521
rect 5342 -572 5362 -148
rect 5426 -572 5446 -148
rect 5874 -199 5978 199
rect 6354 148 6374 572
rect 6438 148 6458 572
rect 6886 521 6990 919
rect 7366 868 7386 1292
rect 7450 868 7470 1292
rect 7366 572 7470 868
rect 6777 520 7099 521
rect 6777 200 6778 520
rect 7098 200 7099 520
rect 6777 199 7099 200
rect 6354 -148 6458 148
rect 5765 -200 6087 -199
rect 5765 -520 5766 -200
rect 6086 -520 6087 -200
rect 5765 -521 6087 -520
rect 5342 -868 5446 -572
rect 4753 -920 5075 -919
rect 4753 -1240 4754 -920
rect 5074 -1240 5075 -920
rect 4753 -1241 5075 -1240
rect 4330 -1588 4434 -1292
rect 3741 -1640 4063 -1639
rect 3741 -1960 3742 -1640
rect 4062 -1960 4063 -1640
rect 3741 -1961 4063 -1960
rect 3318 -2308 3422 -2012
rect 2729 -2360 3051 -2359
rect 2729 -2680 2730 -2360
rect 3050 -2680 3051 -2360
rect 2729 -2681 3051 -2680
rect 2306 -3028 2410 -2732
rect 1717 -3080 2039 -3079
rect 1717 -3400 1718 -3080
rect 2038 -3400 2039 -3080
rect 1717 -3401 2039 -3400
rect 1294 -3748 1398 -3452
rect 705 -3800 1027 -3799
rect 705 -4120 706 -3800
rect 1026 -4120 1027 -3800
rect 705 -4121 1027 -4120
rect 282 -4468 386 -4172
rect -307 -4520 15 -4519
rect -307 -4840 -306 -4520
rect 14 -4840 15 -4520
rect -307 -4841 15 -4840
rect -730 -5188 -626 -4892
rect -1319 -5240 -997 -5239
rect -1319 -5560 -1318 -5240
rect -998 -5560 -997 -5240
rect -1319 -5561 -997 -5560
rect -1742 -5908 -1638 -5612
rect -2331 -5960 -2009 -5959
rect -2331 -6280 -2330 -5960
rect -2010 -6280 -2009 -5960
rect -2331 -6281 -2009 -6280
rect -2754 -6628 -2650 -6332
rect -3343 -6680 -3021 -6679
rect -3343 -7000 -3342 -6680
rect -3022 -7000 -3021 -6680
rect -3343 -7001 -3021 -7000
rect -3766 -7348 -3662 -7052
rect -4355 -7400 -4033 -7399
rect -4355 -7720 -4354 -7400
rect -4034 -7720 -4033 -7400
rect -4355 -7721 -4033 -7720
rect -4778 -8068 -4674 -7772
rect -5367 -8120 -5045 -8119
rect -5367 -8440 -5366 -8120
rect -5046 -8440 -5045 -8120
rect -5367 -8441 -5045 -8440
rect -5790 -8788 -5686 -8492
rect -6379 -8840 -6057 -8839
rect -6379 -9160 -6378 -8840
rect -6058 -9160 -6057 -8840
rect -6379 -9161 -6057 -9160
rect -6802 -9508 -6698 -9212
rect -7391 -9560 -7069 -9559
rect -7391 -9880 -7390 -9560
rect -7070 -9880 -7069 -9560
rect -7391 -9881 -7069 -9880
rect -7282 -10279 -7178 -9881
rect -6802 -9932 -6782 -9508
rect -6718 -9932 -6698 -9508
rect -6270 -9559 -6166 -9161
rect -5790 -9212 -5770 -8788
rect -5706 -9212 -5686 -8788
rect -5258 -8839 -5154 -8441
rect -4778 -8492 -4758 -8068
rect -4694 -8492 -4674 -8068
rect -4246 -8119 -4142 -7721
rect -3766 -7772 -3746 -7348
rect -3682 -7772 -3662 -7348
rect -3234 -7399 -3130 -7001
rect -2754 -7052 -2734 -6628
rect -2670 -7052 -2650 -6628
rect -2222 -6679 -2118 -6281
rect -1742 -6332 -1722 -5908
rect -1658 -6332 -1638 -5908
rect -1210 -5959 -1106 -5561
rect -730 -5612 -710 -5188
rect -646 -5612 -626 -5188
rect -198 -5239 -94 -4841
rect 282 -4892 302 -4468
rect 366 -4892 386 -4468
rect 814 -4519 918 -4121
rect 1294 -4172 1314 -3748
rect 1378 -4172 1398 -3748
rect 1826 -3799 1930 -3401
rect 2306 -3452 2326 -3028
rect 2390 -3452 2410 -3028
rect 2838 -3079 2942 -2681
rect 3318 -2732 3338 -2308
rect 3402 -2732 3422 -2308
rect 3850 -2359 3954 -1961
rect 4330 -2012 4350 -1588
rect 4414 -2012 4434 -1588
rect 4862 -1639 4966 -1241
rect 5342 -1292 5362 -868
rect 5426 -1292 5446 -868
rect 5874 -919 5978 -521
rect 6354 -572 6374 -148
rect 6438 -572 6458 -148
rect 6886 -199 6990 199
rect 7366 148 7386 572
rect 7450 148 7470 572
rect 7366 -148 7470 148
rect 6777 -200 7099 -199
rect 6777 -520 6778 -200
rect 7098 -520 7099 -200
rect 6777 -521 7099 -520
rect 6354 -868 6458 -572
rect 5765 -920 6087 -919
rect 5765 -1240 5766 -920
rect 6086 -1240 6087 -920
rect 5765 -1241 6087 -1240
rect 5342 -1588 5446 -1292
rect 4753 -1640 5075 -1639
rect 4753 -1960 4754 -1640
rect 5074 -1960 5075 -1640
rect 4753 -1961 5075 -1960
rect 4330 -2308 4434 -2012
rect 3741 -2360 4063 -2359
rect 3741 -2680 3742 -2360
rect 4062 -2680 4063 -2360
rect 3741 -2681 4063 -2680
rect 3318 -3028 3422 -2732
rect 2729 -3080 3051 -3079
rect 2729 -3400 2730 -3080
rect 3050 -3400 3051 -3080
rect 2729 -3401 3051 -3400
rect 2306 -3748 2410 -3452
rect 1717 -3800 2039 -3799
rect 1717 -4120 1718 -3800
rect 2038 -4120 2039 -3800
rect 1717 -4121 2039 -4120
rect 1294 -4468 1398 -4172
rect 705 -4520 1027 -4519
rect 705 -4840 706 -4520
rect 1026 -4840 1027 -4520
rect 705 -4841 1027 -4840
rect 282 -5188 386 -4892
rect -307 -5240 15 -5239
rect -307 -5560 -306 -5240
rect 14 -5560 15 -5240
rect -307 -5561 15 -5560
rect -730 -5908 -626 -5612
rect -1319 -5960 -997 -5959
rect -1319 -6280 -1318 -5960
rect -998 -6280 -997 -5960
rect -1319 -6281 -997 -6280
rect -1742 -6628 -1638 -6332
rect -2331 -6680 -2009 -6679
rect -2331 -7000 -2330 -6680
rect -2010 -7000 -2009 -6680
rect -2331 -7001 -2009 -7000
rect -2754 -7348 -2650 -7052
rect -3343 -7400 -3021 -7399
rect -3343 -7720 -3342 -7400
rect -3022 -7720 -3021 -7400
rect -3343 -7721 -3021 -7720
rect -3766 -8068 -3662 -7772
rect -4355 -8120 -4033 -8119
rect -4355 -8440 -4354 -8120
rect -4034 -8440 -4033 -8120
rect -4355 -8441 -4033 -8440
rect -4778 -8788 -4674 -8492
rect -5367 -8840 -5045 -8839
rect -5367 -9160 -5366 -8840
rect -5046 -9160 -5045 -8840
rect -5367 -9161 -5045 -9160
rect -5790 -9508 -5686 -9212
rect -6379 -9560 -6057 -9559
rect -6379 -9880 -6378 -9560
rect -6058 -9880 -6057 -9560
rect -6379 -9881 -6057 -9880
rect -6802 -10228 -6698 -9932
rect -7391 -10280 -7069 -10279
rect -7391 -10600 -7390 -10280
rect -7070 -10600 -7069 -10280
rect -7391 -10601 -7069 -10600
rect -7282 -10999 -7178 -10601
rect -6802 -10652 -6782 -10228
rect -6718 -10652 -6698 -10228
rect -6270 -10279 -6166 -9881
rect -5790 -9932 -5770 -9508
rect -5706 -9932 -5686 -9508
rect -5258 -9559 -5154 -9161
rect -4778 -9212 -4758 -8788
rect -4694 -9212 -4674 -8788
rect -4246 -8839 -4142 -8441
rect -3766 -8492 -3746 -8068
rect -3682 -8492 -3662 -8068
rect -3234 -8119 -3130 -7721
rect -2754 -7772 -2734 -7348
rect -2670 -7772 -2650 -7348
rect -2222 -7399 -2118 -7001
rect -1742 -7052 -1722 -6628
rect -1658 -7052 -1638 -6628
rect -1210 -6679 -1106 -6281
rect -730 -6332 -710 -5908
rect -646 -6332 -626 -5908
rect -198 -5959 -94 -5561
rect 282 -5612 302 -5188
rect 366 -5612 386 -5188
rect 814 -5239 918 -4841
rect 1294 -4892 1314 -4468
rect 1378 -4892 1398 -4468
rect 1826 -4519 1930 -4121
rect 2306 -4172 2326 -3748
rect 2390 -4172 2410 -3748
rect 2838 -3799 2942 -3401
rect 3318 -3452 3338 -3028
rect 3402 -3452 3422 -3028
rect 3850 -3079 3954 -2681
rect 4330 -2732 4350 -2308
rect 4414 -2732 4434 -2308
rect 4862 -2359 4966 -1961
rect 5342 -2012 5362 -1588
rect 5426 -2012 5446 -1588
rect 5874 -1639 5978 -1241
rect 6354 -1292 6374 -868
rect 6438 -1292 6458 -868
rect 6886 -919 6990 -521
rect 7366 -572 7386 -148
rect 7450 -572 7470 -148
rect 7366 -868 7470 -572
rect 6777 -920 7099 -919
rect 6777 -1240 6778 -920
rect 7098 -1240 7099 -920
rect 6777 -1241 7099 -1240
rect 6354 -1588 6458 -1292
rect 5765 -1640 6087 -1639
rect 5765 -1960 5766 -1640
rect 6086 -1960 6087 -1640
rect 5765 -1961 6087 -1960
rect 5342 -2308 5446 -2012
rect 4753 -2360 5075 -2359
rect 4753 -2680 4754 -2360
rect 5074 -2680 5075 -2360
rect 4753 -2681 5075 -2680
rect 4330 -3028 4434 -2732
rect 3741 -3080 4063 -3079
rect 3741 -3400 3742 -3080
rect 4062 -3400 4063 -3080
rect 3741 -3401 4063 -3400
rect 3318 -3748 3422 -3452
rect 2729 -3800 3051 -3799
rect 2729 -4120 2730 -3800
rect 3050 -4120 3051 -3800
rect 2729 -4121 3051 -4120
rect 2306 -4468 2410 -4172
rect 1717 -4520 2039 -4519
rect 1717 -4840 1718 -4520
rect 2038 -4840 2039 -4520
rect 1717 -4841 2039 -4840
rect 1294 -5188 1398 -4892
rect 705 -5240 1027 -5239
rect 705 -5560 706 -5240
rect 1026 -5560 1027 -5240
rect 705 -5561 1027 -5560
rect 282 -5908 386 -5612
rect -307 -5960 15 -5959
rect -307 -6280 -306 -5960
rect 14 -6280 15 -5960
rect -307 -6281 15 -6280
rect -730 -6628 -626 -6332
rect -1319 -6680 -997 -6679
rect -1319 -7000 -1318 -6680
rect -998 -7000 -997 -6680
rect -1319 -7001 -997 -7000
rect -1742 -7348 -1638 -7052
rect -2331 -7400 -2009 -7399
rect -2331 -7720 -2330 -7400
rect -2010 -7720 -2009 -7400
rect -2331 -7721 -2009 -7720
rect -2754 -8068 -2650 -7772
rect -3343 -8120 -3021 -8119
rect -3343 -8440 -3342 -8120
rect -3022 -8440 -3021 -8120
rect -3343 -8441 -3021 -8440
rect -3766 -8788 -3662 -8492
rect -4355 -8840 -4033 -8839
rect -4355 -9160 -4354 -8840
rect -4034 -9160 -4033 -8840
rect -4355 -9161 -4033 -9160
rect -4778 -9508 -4674 -9212
rect -5367 -9560 -5045 -9559
rect -5367 -9880 -5366 -9560
rect -5046 -9880 -5045 -9560
rect -5367 -9881 -5045 -9880
rect -5790 -10228 -5686 -9932
rect -6379 -10280 -6057 -10279
rect -6379 -10600 -6378 -10280
rect -6058 -10600 -6057 -10280
rect -6379 -10601 -6057 -10600
rect -6802 -10948 -6698 -10652
rect -7391 -11000 -7069 -10999
rect -7391 -11320 -7390 -11000
rect -7070 -11320 -7069 -11000
rect -7391 -11321 -7069 -11320
rect -7282 -11520 -7178 -11321
rect -6802 -11372 -6782 -10948
rect -6718 -11372 -6698 -10948
rect -6270 -10999 -6166 -10601
rect -5790 -10652 -5770 -10228
rect -5706 -10652 -5686 -10228
rect -5258 -10279 -5154 -9881
rect -4778 -9932 -4758 -9508
rect -4694 -9932 -4674 -9508
rect -4246 -9559 -4142 -9161
rect -3766 -9212 -3746 -8788
rect -3682 -9212 -3662 -8788
rect -3234 -8839 -3130 -8441
rect -2754 -8492 -2734 -8068
rect -2670 -8492 -2650 -8068
rect -2222 -8119 -2118 -7721
rect -1742 -7772 -1722 -7348
rect -1658 -7772 -1638 -7348
rect -1210 -7399 -1106 -7001
rect -730 -7052 -710 -6628
rect -646 -7052 -626 -6628
rect -198 -6679 -94 -6281
rect 282 -6332 302 -5908
rect 366 -6332 386 -5908
rect 814 -5959 918 -5561
rect 1294 -5612 1314 -5188
rect 1378 -5612 1398 -5188
rect 1826 -5239 1930 -4841
rect 2306 -4892 2326 -4468
rect 2390 -4892 2410 -4468
rect 2838 -4519 2942 -4121
rect 3318 -4172 3338 -3748
rect 3402 -4172 3422 -3748
rect 3850 -3799 3954 -3401
rect 4330 -3452 4350 -3028
rect 4414 -3452 4434 -3028
rect 4862 -3079 4966 -2681
rect 5342 -2732 5362 -2308
rect 5426 -2732 5446 -2308
rect 5874 -2359 5978 -1961
rect 6354 -2012 6374 -1588
rect 6438 -2012 6458 -1588
rect 6886 -1639 6990 -1241
rect 7366 -1292 7386 -868
rect 7450 -1292 7470 -868
rect 7366 -1588 7470 -1292
rect 6777 -1640 7099 -1639
rect 6777 -1960 6778 -1640
rect 7098 -1960 7099 -1640
rect 6777 -1961 7099 -1960
rect 6354 -2308 6458 -2012
rect 5765 -2360 6087 -2359
rect 5765 -2680 5766 -2360
rect 6086 -2680 6087 -2360
rect 5765 -2681 6087 -2680
rect 5342 -3028 5446 -2732
rect 4753 -3080 5075 -3079
rect 4753 -3400 4754 -3080
rect 5074 -3400 5075 -3080
rect 4753 -3401 5075 -3400
rect 4330 -3748 4434 -3452
rect 3741 -3800 4063 -3799
rect 3741 -4120 3742 -3800
rect 4062 -4120 4063 -3800
rect 3741 -4121 4063 -4120
rect 3318 -4468 3422 -4172
rect 2729 -4520 3051 -4519
rect 2729 -4840 2730 -4520
rect 3050 -4840 3051 -4520
rect 2729 -4841 3051 -4840
rect 2306 -5188 2410 -4892
rect 1717 -5240 2039 -5239
rect 1717 -5560 1718 -5240
rect 2038 -5560 2039 -5240
rect 1717 -5561 2039 -5560
rect 1294 -5908 1398 -5612
rect 705 -5960 1027 -5959
rect 705 -6280 706 -5960
rect 1026 -6280 1027 -5960
rect 705 -6281 1027 -6280
rect 282 -6628 386 -6332
rect -307 -6680 15 -6679
rect -307 -7000 -306 -6680
rect 14 -7000 15 -6680
rect -307 -7001 15 -7000
rect -730 -7348 -626 -7052
rect -1319 -7400 -997 -7399
rect -1319 -7720 -1318 -7400
rect -998 -7720 -997 -7400
rect -1319 -7721 -997 -7720
rect -1742 -8068 -1638 -7772
rect -2331 -8120 -2009 -8119
rect -2331 -8440 -2330 -8120
rect -2010 -8440 -2009 -8120
rect -2331 -8441 -2009 -8440
rect -2754 -8788 -2650 -8492
rect -3343 -8840 -3021 -8839
rect -3343 -9160 -3342 -8840
rect -3022 -9160 -3021 -8840
rect -3343 -9161 -3021 -9160
rect -3766 -9508 -3662 -9212
rect -4355 -9560 -4033 -9559
rect -4355 -9880 -4354 -9560
rect -4034 -9880 -4033 -9560
rect -4355 -9881 -4033 -9880
rect -4778 -10228 -4674 -9932
rect -5367 -10280 -5045 -10279
rect -5367 -10600 -5366 -10280
rect -5046 -10600 -5045 -10280
rect -5367 -10601 -5045 -10600
rect -5790 -10948 -5686 -10652
rect -6379 -11000 -6057 -10999
rect -6379 -11320 -6378 -11000
rect -6058 -11320 -6057 -11000
rect -6379 -11321 -6057 -11320
rect -6802 -11520 -6698 -11372
rect -6270 -11520 -6166 -11321
rect -5790 -11372 -5770 -10948
rect -5706 -11372 -5686 -10948
rect -5258 -10999 -5154 -10601
rect -4778 -10652 -4758 -10228
rect -4694 -10652 -4674 -10228
rect -4246 -10279 -4142 -9881
rect -3766 -9932 -3746 -9508
rect -3682 -9932 -3662 -9508
rect -3234 -9559 -3130 -9161
rect -2754 -9212 -2734 -8788
rect -2670 -9212 -2650 -8788
rect -2222 -8839 -2118 -8441
rect -1742 -8492 -1722 -8068
rect -1658 -8492 -1638 -8068
rect -1210 -8119 -1106 -7721
rect -730 -7772 -710 -7348
rect -646 -7772 -626 -7348
rect -198 -7399 -94 -7001
rect 282 -7052 302 -6628
rect 366 -7052 386 -6628
rect 814 -6679 918 -6281
rect 1294 -6332 1314 -5908
rect 1378 -6332 1398 -5908
rect 1826 -5959 1930 -5561
rect 2306 -5612 2326 -5188
rect 2390 -5612 2410 -5188
rect 2838 -5239 2942 -4841
rect 3318 -4892 3338 -4468
rect 3402 -4892 3422 -4468
rect 3850 -4519 3954 -4121
rect 4330 -4172 4350 -3748
rect 4414 -4172 4434 -3748
rect 4862 -3799 4966 -3401
rect 5342 -3452 5362 -3028
rect 5426 -3452 5446 -3028
rect 5874 -3079 5978 -2681
rect 6354 -2732 6374 -2308
rect 6438 -2732 6458 -2308
rect 6886 -2359 6990 -1961
rect 7366 -2012 7386 -1588
rect 7450 -2012 7470 -1588
rect 7366 -2308 7470 -2012
rect 6777 -2360 7099 -2359
rect 6777 -2680 6778 -2360
rect 7098 -2680 7099 -2360
rect 6777 -2681 7099 -2680
rect 6354 -3028 6458 -2732
rect 5765 -3080 6087 -3079
rect 5765 -3400 5766 -3080
rect 6086 -3400 6087 -3080
rect 5765 -3401 6087 -3400
rect 5342 -3748 5446 -3452
rect 4753 -3800 5075 -3799
rect 4753 -4120 4754 -3800
rect 5074 -4120 5075 -3800
rect 4753 -4121 5075 -4120
rect 4330 -4468 4434 -4172
rect 3741 -4520 4063 -4519
rect 3741 -4840 3742 -4520
rect 4062 -4840 4063 -4520
rect 3741 -4841 4063 -4840
rect 3318 -5188 3422 -4892
rect 2729 -5240 3051 -5239
rect 2729 -5560 2730 -5240
rect 3050 -5560 3051 -5240
rect 2729 -5561 3051 -5560
rect 2306 -5908 2410 -5612
rect 1717 -5960 2039 -5959
rect 1717 -6280 1718 -5960
rect 2038 -6280 2039 -5960
rect 1717 -6281 2039 -6280
rect 1294 -6628 1398 -6332
rect 705 -6680 1027 -6679
rect 705 -7000 706 -6680
rect 1026 -7000 1027 -6680
rect 705 -7001 1027 -7000
rect 282 -7348 386 -7052
rect -307 -7400 15 -7399
rect -307 -7720 -306 -7400
rect 14 -7720 15 -7400
rect -307 -7721 15 -7720
rect -730 -8068 -626 -7772
rect -1319 -8120 -997 -8119
rect -1319 -8440 -1318 -8120
rect -998 -8440 -997 -8120
rect -1319 -8441 -997 -8440
rect -1742 -8788 -1638 -8492
rect -2331 -8840 -2009 -8839
rect -2331 -9160 -2330 -8840
rect -2010 -9160 -2009 -8840
rect -2331 -9161 -2009 -9160
rect -2754 -9508 -2650 -9212
rect -3343 -9560 -3021 -9559
rect -3343 -9880 -3342 -9560
rect -3022 -9880 -3021 -9560
rect -3343 -9881 -3021 -9880
rect -3766 -10228 -3662 -9932
rect -4355 -10280 -4033 -10279
rect -4355 -10600 -4354 -10280
rect -4034 -10600 -4033 -10280
rect -4355 -10601 -4033 -10600
rect -4778 -10948 -4674 -10652
rect -5367 -11000 -5045 -10999
rect -5367 -11320 -5366 -11000
rect -5046 -11320 -5045 -11000
rect -5367 -11321 -5045 -11320
rect -5790 -11520 -5686 -11372
rect -5258 -11520 -5154 -11321
rect -4778 -11372 -4758 -10948
rect -4694 -11372 -4674 -10948
rect -4246 -10999 -4142 -10601
rect -3766 -10652 -3746 -10228
rect -3682 -10652 -3662 -10228
rect -3234 -10279 -3130 -9881
rect -2754 -9932 -2734 -9508
rect -2670 -9932 -2650 -9508
rect -2222 -9559 -2118 -9161
rect -1742 -9212 -1722 -8788
rect -1658 -9212 -1638 -8788
rect -1210 -8839 -1106 -8441
rect -730 -8492 -710 -8068
rect -646 -8492 -626 -8068
rect -198 -8119 -94 -7721
rect 282 -7772 302 -7348
rect 366 -7772 386 -7348
rect 814 -7399 918 -7001
rect 1294 -7052 1314 -6628
rect 1378 -7052 1398 -6628
rect 1826 -6679 1930 -6281
rect 2306 -6332 2326 -5908
rect 2390 -6332 2410 -5908
rect 2838 -5959 2942 -5561
rect 3318 -5612 3338 -5188
rect 3402 -5612 3422 -5188
rect 3850 -5239 3954 -4841
rect 4330 -4892 4350 -4468
rect 4414 -4892 4434 -4468
rect 4862 -4519 4966 -4121
rect 5342 -4172 5362 -3748
rect 5426 -4172 5446 -3748
rect 5874 -3799 5978 -3401
rect 6354 -3452 6374 -3028
rect 6438 -3452 6458 -3028
rect 6886 -3079 6990 -2681
rect 7366 -2732 7386 -2308
rect 7450 -2732 7470 -2308
rect 7366 -3028 7470 -2732
rect 6777 -3080 7099 -3079
rect 6777 -3400 6778 -3080
rect 7098 -3400 7099 -3080
rect 6777 -3401 7099 -3400
rect 6354 -3748 6458 -3452
rect 5765 -3800 6087 -3799
rect 5765 -4120 5766 -3800
rect 6086 -4120 6087 -3800
rect 5765 -4121 6087 -4120
rect 5342 -4468 5446 -4172
rect 4753 -4520 5075 -4519
rect 4753 -4840 4754 -4520
rect 5074 -4840 5075 -4520
rect 4753 -4841 5075 -4840
rect 4330 -5188 4434 -4892
rect 3741 -5240 4063 -5239
rect 3741 -5560 3742 -5240
rect 4062 -5560 4063 -5240
rect 3741 -5561 4063 -5560
rect 3318 -5908 3422 -5612
rect 2729 -5960 3051 -5959
rect 2729 -6280 2730 -5960
rect 3050 -6280 3051 -5960
rect 2729 -6281 3051 -6280
rect 2306 -6628 2410 -6332
rect 1717 -6680 2039 -6679
rect 1717 -7000 1718 -6680
rect 2038 -7000 2039 -6680
rect 1717 -7001 2039 -7000
rect 1294 -7348 1398 -7052
rect 705 -7400 1027 -7399
rect 705 -7720 706 -7400
rect 1026 -7720 1027 -7400
rect 705 -7721 1027 -7720
rect 282 -8068 386 -7772
rect -307 -8120 15 -8119
rect -307 -8440 -306 -8120
rect 14 -8440 15 -8120
rect -307 -8441 15 -8440
rect -730 -8788 -626 -8492
rect -1319 -8840 -997 -8839
rect -1319 -9160 -1318 -8840
rect -998 -9160 -997 -8840
rect -1319 -9161 -997 -9160
rect -1742 -9508 -1638 -9212
rect -2331 -9560 -2009 -9559
rect -2331 -9880 -2330 -9560
rect -2010 -9880 -2009 -9560
rect -2331 -9881 -2009 -9880
rect -2754 -10228 -2650 -9932
rect -3343 -10280 -3021 -10279
rect -3343 -10600 -3342 -10280
rect -3022 -10600 -3021 -10280
rect -3343 -10601 -3021 -10600
rect -3766 -10948 -3662 -10652
rect -4355 -11000 -4033 -10999
rect -4355 -11320 -4354 -11000
rect -4034 -11320 -4033 -11000
rect -4355 -11321 -4033 -11320
rect -4778 -11520 -4674 -11372
rect -4246 -11520 -4142 -11321
rect -3766 -11372 -3746 -10948
rect -3682 -11372 -3662 -10948
rect -3234 -10999 -3130 -10601
rect -2754 -10652 -2734 -10228
rect -2670 -10652 -2650 -10228
rect -2222 -10279 -2118 -9881
rect -1742 -9932 -1722 -9508
rect -1658 -9932 -1638 -9508
rect -1210 -9559 -1106 -9161
rect -730 -9212 -710 -8788
rect -646 -9212 -626 -8788
rect -198 -8839 -94 -8441
rect 282 -8492 302 -8068
rect 366 -8492 386 -8068
rect 814 -8119 918 -7721
rect 1294 -7772 1314 -7348
rect 1378 -7772 1398 -7348
rect 1826 -7399 1930 -7001
rect 2306 -7052 2326 -6628
rect 2390 -7052 2410 -6628
rect 2838 -6679 2942 -6281
rect 3318 -6332 3338 -5908
rect 3402 -6332 3422 -5908
rect 3850 -5959 3954 -5561
rect 4330 -5612 4350 -5188
rect 4414 -5612 4434 -5188
rect 4862 -5239 4966 -4841
rect 5342 -4892 5362 -4468
rect 5426 -4892 5446 -4468
rect 5874 -4519 5978 -4121
rect 6354 -4172 6374 -3748
rect 6438 -4172 6458 -3748
rect 6886 -3799 6990 -3401
rect 7366 -3452 7386 -3028
rect 7450 -3452 7470 -3028
rect 7366 -3748 7470 -3452
rect 6777 -3800 7099 -3799
rect 6777 -4120 6778 -3800
rect 7098 -4120 7099 -3800
rect 6777 -4121 7099 -4120
rect 6354 -4468 6458 -4172
rect 5765 -4520 6087 -4519
rect 5765 -4840 5766 -4520
rect 6086 -4840 6087 -4520
rect 5765 -4841 6087 -4840
rect 5342 -5188 5446 -4892
rect 4753 -5240 5075 -5239
rect 4753 -5560 4754 -5240
rect 5074 -5560 5075 -5240
rect 4753 -5561 5075 -5560
rect 4330 -5908 4434 -5612
rect 3741 -5960 4063 -5959
rect 3741 -6280 3742 -5960
rect 4062 -6280 4063 -5960
rect 3741 -6281 4063 -6280
rect 3318 -6628 3422 -6332
rect 2729 -6680 3051 -6679
rect 2729 -7000 2730 -6680
rect 3050 -7000 3051 -6680
rect 2729 -7001 3051 -7000
rect 2306 -7348 2410 -7052
rect 1717 -7400 2039 -7399
rect 1717 -7720 1718 -7400
rect 2038 -7720 2039 -7400
rect 1717 -7721 2039 -7720
rect 1294 -8068 1398 -7772
rect 705 -8120 1027 -8119
rect 705 -8440 706 -8120
rect 1026 -8440 1027 -8120
rect 705 -8441 1027 -8440
rect 282 -8788 386 -8492
rect -307 -8840 15 -8839
rect -307 -9160 -306 -8840
rect 14 -9160 15 -8840
rect -307 -9161 15 -9160
rect -730 -9508 -626 -9212
rect -1319 -9560 -997 -9559
rect -1319 -9880 -1318 -9560
rect -998 -9880 -997 -9560
rect -1319 -9881 -997 -9880
rect -1742 -10228 -1638 -9932
rect -2331 -10280 -2009 -10279
rect -2331 -10600 -2330 -10280
rect -2010 -10600 -2009 -10280
rect -2331 -10601 -2009 -10600
rect -2754 -10948 -2650 -10652
rect -3343 -11000 -3021 -10999
rect -3343 -11320 -3342 -11000
rect -3022 -11320 -3021 -11000
rect -3343 -11321 -3021 -11320
rect -3766 -11520 -3662 -11372
rect -3234 -11520 -3130 -11321
rect -2754 -11372 -2734 -10948
rect -2670 -11372 -2650 -10948
rect -2222 -10999 -2118 -10601
rect -1742 -10652 -1722 -10228
rect -1658 -10652 -1638 -10228
rect -1210 -10279 -1106 -9881
rect -730 -9932 -710 -9508
rect -646 -9932 -626 -9508
rect -198 -9559 -94 -9161
rect 282 -9212 302 -8788
rect 366 -9212 386 -8788
rect 814 -8839 918 -8441
rect 1294 -8492 1314 -8068
rect 1378 -8492 1398 -8068
rect 1826 -8119 1930 -7721
rect 2306 -7772 2326 -7348
rect 2390 -7772 2410 -7348
rect 2838 -7399 2942 -7001
rect 3318 -7052 3338 -6628
rect 3402 -7052 3422 -6628
rect 3850 -6679 3954 -6281
rect 4330 -6332 4350 -5908
rect 4414 -6332 4434 -5908
rect 4862 -5959 4966 -5561
rect 5342 -5612 5362 -5188
rect 5426 -5612 5446 -5188
rect 5874 -5239 5978 -4841
rect 6354 -4892 6374 -4468
rect 6438 -4892 6458 -4468
rect 6886 -4519 6990 -4121
rect 7366 -4172 7386 -3748
rect 7450 -4172 7470 -3748
rect 7366 -4468 7470 -4172
rect 6777 -4520 7099 -4519
rect 6777 -4840 6778 -4520
rect 7098 -4840 7099 -4520
rect 6777 -4841 7099 -4840
rect 6354 -5188 6458 -4892
rect 5765 -5240 6087 -5239
rect 5765 -5560 5766 -5240
rect 6086 -5560 6087 -5240
rect 5765 -5561 6087 -5560
rect 5342 -5908 5446 -5612
rect 4753 -5960 5075 -5959
rect 4753 -6280 4754 -5960
rect 5074 -6280 5075 -5960
rect 4753 -6281 5075 -6280
rect 4330 -6628 4434 -6332
rect 3741 -6680 4063 -6679
rect 3741 -7000 3742 -6680
rect 4062 -7000 4063 -6680
rect 3741 -7001 4063 -7000
rect 3318 -7348 3422 -7052
rect 2729 -7400 3051 -7399
rect 2729 -7720 2730 -7400
rect 3050 -7720 3051 -7400
rect 2729 -7721 3051 -7720
rect 2306 -8068 2410 -7772
rect 1717 -8120 2039 -8119
rect 1717 -8440 1718 -8120
rect 2038 -8440 2039 -8120
rect 1717 -8441 2039 -8440
rect 1294 -8788 1398 -8492
rect 705 -8840 1027 -8839
rect 705 -9160 706 -8840
rect 1026 -9160 1027 -8840
rect 705 -9161 1027 -9160
rect 282 -9508 386 -9212
rect -307 -9560 15 -9559
rect -307 -9880 -306 -9560
rect 14 -9880 15 -9560
rect -307 -9881 15 -9880
rect -730 -10228 -626 -9932
rect -1319 -10280 -997 -10279
rect -1319 -10600 -1318 -10280
rect -998 -10600 -997 -10280
rect -1319 -10601 -997 -10600
rect -1742 -10948 -1638 -10652
rect -2331 -11000 -2009 -10999
rect -2331 -11320 -2330 -11000
rect -2010 -11320 -2009 -11000
rect -2331 -11321 -2009 -11320
rect -2754 -11520 -2650 -11372
rect -2222 -11520 -2118 -11321
rect -1742 -11372 -1722 -10948
rect -1658 -11372 -1638 -10948
rect -1210 -10999 -1106 -10601
rect -730 -10652 -710 -10228
rect -646 -10652 -626 -10228
rect -198 -10279 -94 -9881
rect 282 -9932 302 -9508
rect 366 -9932 386 -9508
rect 814 -9559 918 -9161
rect 1294 -9212 1314 -8788
rect 1378 -9212 1398 -8788
rect 1826 -8839 1930 -8441
rect 2306 -8492 2326 -8068
rect 2390 -8492 2410 -8068
rect 2838 -8119 2942 -7721
rect 3318 -7772 3338 -7348
rect 3402 -7772 3422 -7348
rect 3850 -7399 3954 -7001
rect 4330 -7052 4350 -6628
rect 4414 -7052 4434 -6628
rect 4862 -6679 4966 -6281
rect 5342 -6332 5362 -5908
rect 5426 -6332 5446 -5908
rect 5874 -5959 5978 -5561
rect 6354 -5612 6374 -5188
rect 6438 -5612 6458 -5188
rect 6886 -5239 6990 -4841
rect 7366 -4892 7386 -4468
rect 7450 -4892 7470 -4468
rect 7366 -5188 7470 -4892
rect 6777 -5240 7099 -5239
rect 6777 -5560 6778 -5240
rect 7098 -5560 7099 -5240
rect 6777 -5561 7099 -5560
rect 6354 -5908 6458 -5612
rect 5765 -5960 6087 -5959
rect 5765 -6280 5766 -5960
rect 6086 -6280 6087 -5960
rect 5765 -6281 6087 -6280
rect 5342 -6628 5446 -6332
rect 4753 -6680 5075 -6679
rect 4753 -7000 4754 -6680
rect 5074 -7000 5075 -6680
rect 4753 -7001 5075 -7000
rect 4330 -7348 4434 -7052
rect 3741 -7400 4063 -7399
rect 3741 -7720 3742 -7400
rect 4062 -7720 4063 -7400
rect 3741 -7721 4063 -7720
rect 3318 -8068 3422 -7772
rect 2729 -8120 3051 -8119
rect 2729 -8440 2730 -8120
rect 3050 -8440 3051 -8120
rect 2729 -8441 3051 -8440
rect 2306 -8788 2410 -8492
rect 1717 -8840 2039 -8839
rect 1717 -9160 1718 -8840
rect 2038 -9160 2039 -8840
rect 1717 -9161 2039 -9160
rect 1294 -9508 1398 -9212
rect 705 -9560 1027 -9559
rect 705 -9880 706 -9560
rect 1026 -9880 1027 -9560
rect 705 -9881 1027 -9880
rect 282 -10228 386 -9932
rect -307 -10280 15 -10279
rect -307 -10600 -306 -10280
rect 14 -10600 15 -10280
rect -307 -10601 15 -10600
rect -730 -10948 -626 -10652
rect -1319 -11000 -997 -10999
rect -1319 -11320 -1318 -11000
rect -998 -11320 -997 -11000
rect -1319 -11321 -997 -11320
rect -1742 -11520 -1638 -11372
rect -1210 -11520 -1106 -11321
rect -730 -11372 -710 -10948
rect -646 -11372 -626 -10948
rect -198 -10999 -94 -10601
rect 282 -10652 302 -10228
rect 366 -10652 386 -10228
rect 814 -10279 918 -9881
rect 1294 -9932 1314 -9508
rect 1378 -9932 1398 -9508
rect 1826 -9559 1930 -9161
rect 2306 -9212 2326 -8788
rect 2390 -9212 2410 -8788
rect 2838 -8839 2942 -8441
rect 3318 -8492 3338 -8068
rect 3402 -8492 3422 -8068
rect 3850 -8119 3954 -7721
rect 4330 -7772 4350 -7348
rect 4414 -7772 4434 -7348
rect 4862 -7399 4966 -7001
rect 5342 -7052 5362 -6628
rect 5426 -7052 5446 -6628
rect 5874 -6679 5978 -6281
rect 6354 -6332 6374 -5908
rect 6438 -6332 6458 -5908
rect 6886 -5959 6990 -5561
rect 7366 -5612 7386 -5188
rect 7450 -5612 7470 -5188
rect 7366 -5908 7470 -5612
rect 6777 -5960 7099 -5959
rect 6777 -6280 6778 -5960
rect 7098 -6280 7099 -5960
rect 6777 -6281 7099 -6280
rect 6354 -6628 6458 -6332
rect 5765 -6680 6087 -6679
rect 5765 -7000 5766 -6680
rect 6086 -7000 6087 -6680
rect 5765 -7001 6087 -7000
rect 5342 -7348 5446 -7052
rect 4753 -7400 5075 -7399
rect 4753 -7720 4754 -7400
rect 5074 -7720 5075 -7400
rect 4753 -7721 5075 -7720
rect 4330 -8068 4434 -7772
rect 3741 -8120 4063 -8119
rect 3741 -8440 3742 -8120
rect 4062 -8440 4063 -8120
rect 3741 -8441 4063 -8440
rect 3318 -8788 3422 -8492
rect 2729 -8840 3051 -8839
rect 2729 -9160 2730 -8840
rect 3050 -9160 3051 -8840
rect 2729 -9161 3051 -9160
rect 2306 -9508 2410 -9212
rect 1717 -9560 2039 -9559
rect 1717 -9880 1718 -9560
rect 2038 -9880 2039 -9560
rect 1717 -9881 2039 -9880
rect 1294 -10228 1398 -9932
rect 705 -10280 1027 -10279
rect 705 -10600 706 -10280
rect 1026 -10600 1027 -10280
rect 705 -10601 1027 -10600
rect 282 -10948 386 -10652
rect -307 -11000 15 -10999
rect -307 -11320 -306 -11000
rect 14 -11320 15 -11000
rect -307 -11321 15 -11320
rect -730 -11520 -626 -11372
rect -198 -11520 -94 -11321
rect 282 -11372 302 -10948
rect 366 -11372 386 -10948
rect 814 -10999 918 -10601
rect 1294 -10652 1314 -10228
rect 1378 -10652 1398 -10228
rect 1826 -10279 1930 -9881
rect 2306 -9932 2326 -9508
rect 2390 -9932 2410 -9508
rect 2838 -9559 2942 -9161
rect 3318 -9212 3338 -8788
rect 3402 -9212 3422 -8788
rect 3850 -8839 3954 -8441
rect 4330 -8492 4350 -8068
rect 4414 -8492 4434 -8068
rect 4862 -8119 4966 -7721
rect 5342 -7772 5362 -7348
rect 5426 -7772 5446 -7348
rect 5874 -7399 5978 -7001
rect 6354 -7052 6374 -6628
rect 6438 -7052 6458 -6628
rect 6886 -6679 6990 -6281
rect 7366 -6332 7386 -5908
rect 7450 -6332 7470 -5908
rect 7366 -6628 7470 -6332
rect 6777 -6680 7099 -6679
rect 6777 -7000 6778 -6680
rect 7098 -7000 7099 -6680
rect 6777 -7001 7099 -7000
rect 6354 -7348 6458 -7052
rect 5765 -7400 6087 -7399
rect 5765 -7720 5766 -7400
rect 6086 -7720 6087 -7400
rect 5765 -7721 6087 -7720
rect 5342 -8068 5446 -7772
rect 4753 -8120 5075 -8119
rect 4753 -8440 4754 -8120
rect 5074 -8440 5075 -8120
rect 4753 -8441 5075 -8440
rect 4330 -8788 4434 -8492
rect 3741 -8840 4063 -8839
rect 3741 -9160 3742 -8840
rect 4062 -9160 4063 -8840
rect 3741 -9161 4063 -9160
rect 3318 -9508 3422 -9212
rect 2729 -9560 3051 -9559
rect 2729 -9880 2730 -9560
rect 3050 -9880 3051 -9560
rect 2729 -9881 3051 -9880
rect 2306 -10228 2410 -9932
rect 1717 -10280 2039 -10279
rect 1717 -10600 1718 -10280
rect 2038 -10600 2039 -10280
rect 1717 -10601 2039 -10600
rect 1294 -10948 1398 -10652
rect 705 -11000 1027 -10999
rect 705 -11320 706 -11000
rect 1026 -11320 1027 -11000
rect 705 -11321 1027 -11320
rect 282 -11520 386 -11372
rect 814 -11520 918 -11321
rect 1294 -11372 1314 -10948
rect 1378 -11372 1398 -10948
rect 1826 -10999 1930 -10601
rect 2306 -10652 2326 -10228
rect 2390 -10652 2410 -10228
rect 2838 -10279 2942 -9881
rect 3318 -9932 3338 -9508
rect 3402 -9932 3422 -9508
rect 3850 -9559 3954 -9161
rect 4330 -9212 4350 -8788
rect 4414 -9212 4434 -8788
rect 4862 -8839 4966 -8441
rect 5342 -8492 5362 -8068
rect 5426 -8492 5446 -8068
rect 5874 -8119 5978 -7721
rect 6354 -7772 6374 -7348
rect 6438 -7772 6458 -7348
rect 6886 -7399 6990 -7001
rect 7366 -7052 7386 -6628
rect 7450 -7052 7470 -6628
rect 7366 -7348 7470 -7052
rect 6777 -7400 7099 -7399
rect 6777 -7720 6778 -7400
rect 7098 -7720 7099 -7400
rect 6777 -7721 7099 -7720
rect 6354 -8068 6458 -7772
rect 5765 -8120 6087 -8119
rect 5765 -8440 5766 -8120
rect 6086 -8440 6087 -8120
rect 5765 -8441 6087 -8440
rect 5342 -8788 5446 -8492
rect 4753 -8840 5075 -8839
rect 4753 -9160 4754 -8840
rect 5074 -9160 5075 -8840
rect 4753 -9161 5075 -9160
rect 4330 -9508 4434 -9212
rect 3741 -9560 4063 -9559
rect 3741 -9880 3742 -9560
rect 4062 -9880 4063 -9560
rect 3741 -9881 4063 -9880
rect 3318 -10228 3422 -9932
rect 2729 -10280 3051 -10279
rect 2729 -10600 2730 -10280
rect 3050 -10600 3051 -10280
rect 2729 -10601 3051 -10600
rect 2306 -10948 2410 -10652
rect 1717 -11000 2039 -10999
rect 1717 -11320 1718 -11000
rect 2038 -11320 2039 -11000
rect 1717 -11321 2039 -11320
rect 1294 -11520 1398 -11372
rect 1826 -11520 1930 -11321
rect 2306 -11372 2326 -10948
rect 2390 -11372 2410 -10948
rect 2838 -10999 2942 -10601
rect 3318 -10652 3338 -10228
rect 3402 -10652 3422 -10228
rect 3850 -10279 3954 -9881
rect 4330 -9932 4350 -9508
rect 4414 -9932 4434 -9508
rect 4862 -9559 4966 -9161
rect 5342 -9212 5362 -8788
rect 5426 -9212 5446 -8788
rect 5874 -8839 5978 -8441
rect 6354 -8492 6374 -8068
rect 6438 -8492 6458 -8068
rect 6886 -8119 6990 -7721
rect 7366 -7772 7386 -7348
rect 7450 -7772 7470 -7348
rect 7366 -8068 7470 -7772
rect 6777 -8120 7099 -8119
rect 6777 -8440 6778 -8120
rect 7098 -8440 7099 -8120
rect 6777 -8441 7099 -8440
rect 6354 -8788 6458 -8492
rect 5765 -8840 6087 -8839
rect 5765 -9160 5766 -8840
rect 6086 -9160 6087 -8840
rect 5765 -9161 6087 -9160
rect 5342 -9508 5446 -9212
rect 4753 -9560 5075 -9559
rect 4753 -9880 4754 -9560
rect 5074 -9880 5075 -9560
rect 4753 -9881 5075 -9880
rect 4330 -10228 4434 -9932
rect 3741 -10280 4063 -10279
rect 3741 -10600 3742 -10280
rect 4062 -10600 4063 -10280
rect 3741 -10601 4063 -10600
rect 3318 -10948 3422 -10652
rect 2729 -11000 3051 -10999
rect 2729 -11320 2730 -11000
rect 3050 -11320 3051 -11000
rect 2729 -11321 3051 -11320
rect 2306 -11520 2410 -11372
rect 2838 -11520 2942 -11321
rect 3318 -11372 3338 -10948
rect 3402 -11372 3422 -10948
rect 3850 -10999 3954 -10601
rect 4330 -10652 4350 -10228
rect 4414 -10652 4434 -10228
rect 4862 -10279 4966 -9881
rect 5342 -9932 5362 -9508
rect 5426 -9932 5446 -9508
rect 5874 -9559 5978 -9161
rect 6354 -9212 6374 -8788
rect 6438 -9212 6458 -8788
rect 6886 -8839 6990 -8441
rect 7366 -8492 7386 -8068
rect 7450 -8492 7470 -8068
rect 7366 -8788 7470 -8492
rect 6777 -8840 7099 -8839
rect 6777 -9160 6778 -8840
rect 7098 -9160 7099 -8840
rect 6777 -9161 7099 -9160
rect 6354 -9508 6458 -9212
rect 5765 -9560 6087 -9559
rect 5765 -9880 5766 -9560
rect 6086 -9880 6087 -9560
rect 5765 -9881 6087 -9880
rect 5342 -10228 5446 -9932
rect 4753 -10280 5075 -10279
rect 4753 -10600 4754 -10280
rect 5074 -10600 5075 -10280
rect 4753 -10601 5075 -10600
rect 4330 -10948 4434 -10652
rect 3741 -11000 4063 -10999
rect 3741 -11320 3742 -11000
rect 4062 -11320 4063 -11000
rect 3741 -11321 4063 -11320
rect 3318 -11520 3422 -11372
rect 3850 -11520 3954 -11321
rect 4330 -11372 4350 -10948
rect 4414 -11372 4434 -10948
rect 4862 -10999 4966 -10601
rect 5342 -10652 5362 -10228
rect 5426 -10652 5446 -10228
rect 5874 -10279 5978 -9881
rect 6354 -9932 6374 -9508
rect 6438 -9932 6458 -9508
rect 6886 -9559 6990 -9161
rect 7366 -9212 7386 -8788
rect 7450 -9212 7470 -8788
rect 7366 -9508 7470 -9212
rect 6777 -9560 7099 -9559
rect 6777 -9880 6778 -9560
rect 7098 -9880 7099 -9560
rect 6777 -9881 7099 -9880
rect 6354 -10228 6458 -9932
rect 5765 -10280 6087 -10279
rect 5765 -10600 5766 -10280
rect 6086 -10600 6087 -10280
rect 5765 -10601 6087 -10600
rect 5342 -10948 5446 -10652
rect 4753 -11000 5075 -10999
rect 4753 -11320 4754 -11000
rect 5074 -11320 5075 -11000
rect 4753 -11321 5075 -11320
rect 4330 -11520 4434 -11372
rect 4862 -11520 4966 -11321
rect 5342 -11372 5362 -10948
rect 5426 -11372 5446 -10948
rect 5874 -10999 5978 -10601
rect 6354 -10652 6374 -10228
rect 6438 -10652 6458 -10228
rect 6886 -10279 6990 -9881
rect 7366 -9932 7386 -9508
rect 7450 -9932 7470 -9508
rect 7366 -10228 7470 -9932
rect 6777 -10280 7099 -10279
rect 6777 -10600 6778 -10280
rect 7098 -10600 7099 -10280
rect 6777 -10601 7099 -10600
rect 6354 -10948 6458 -10652
rect 5765 -11000 6087 -10999
rect 5765 -11320 5766 -11000
rect 6086 -11320 6087 -11000
rect 5765 -11321 6087 -11320
rect 5342 -11520 5446 -11372
rect 5874 -11520 5978 -11321
rect 6354 -11372 6374 -10948
rect 6438 -11372 6458 -10948
rect 6886 -10999 6990 -10601
rect 7366 -10652 7386 -10228
rect 7450 -10652 7470 -10228
rect 7366 -10948 7470 -10652
rect 6777 -11000 7099 -10999
rect 6777 -11320 6778 -11000
rect 7098 -11320 7099 -11000
rect 6777 -11321 7099 -11320
rect 6354 -11520 6458 -11372
rect 6886 -11520 6990 -11321
rect 7366 -11372 7386 -10948
rect 7450 -11372 7470 -10948
rect 7366 -11520 7470 -11372
<< properties >>
string FIXED_BBOX 6698 10920 7178 11400
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 15 ny 32 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
