magic
tech sky130A
magscale 1 2
timestamp 1729087186
<< error_p >>
rect -29 541 29 547
rect -29 507 -17 541
rect -29 501 29 507
<< pwell >>
rect -226 -679 226 679
<< nmos >>
rect -30 -531 30 469
<< ndiff >>
rect -88 457 -30 469
rect -88 -519 -76 457
rect -42 -519 -30 457
rect -88 -531 -30 -519
rect 30 457 88 469
rect 30 -519 42 457
rect 76 -519 88 457
rect 30 -531 88 -519
<< ndiffc >>
rect -76 -519 -42 457
rect 42 -519 76 457
<< psubdiff >>
rect -190 609 -94 643
rect 94 609 190 643
rect -190 547 -156 609
rect 156 547 190 609
rect -190 -609 -156 -547
rect 156 -609 190 -547
rect -190 -643 -94 -609
rect 94 -643 190 -609
<< psubdiffcont >>
rect -94 609 94 643
rect -190 -547 -156 547
rect 156 -547 190 547
rect -94 -643 94 -609
<< poly >>
rect -33 541 33 557
rect -33 507 -17 541
rect 17 507 33 541
rect -33 491 33 507
rect -30 469 30 491
rect -30 -557 30 -531
<< polycont >>
rect -17 507 17 541
<< locali >>
rect -190 609 -94 643
rect 94 609 190 643
rect -190 547 -156 609
rect 156 547 190 609
rect -33 507 -17 541
rect 17 507 33 541
rect -76 457 -42 473
rect -76 -535 -42 -519
rect 42 457 76 473
rect 42 -535 76 -519
rect -190 -609 -156 -547
rect 156 -609 190 -547
rect -190 -643 -94 -609
rect 94 -643 190 -609
<< viali >>
rect -17 507 17 541
rect -76 -519 -42 457
rect 42 -519 76 457
<< metal1 >>
rect -29 541 29 547
rect -29 507 -17 541
rect 17 507 29 541
rect -29 501 29 507
rect -82 457 -36 469
rect -82 -519 -76 457
rect -42 -519 -36 457
rect -82 -531 -36 -519
rect 36 457 82 469
rect 36 -519 42 457
rect 76 -519 82 457
rect 36 -531 82 -519
<< properties >>
string FIXED_BBOX -173 -626 173 626
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
