magic
tech sky130A
magscale 1 2
timestamp 1730624594
<< nwell >>
rect -246 -637 246 637
<< pmos >>
rect -50 118 50 418
rect -50 -418 50 -118
<< pdiff >>
rect -108 406 -50 418
rect -108 130 -96 406
rect -62 130 -50 406
rect -108 118 -50 130
rect 50 406 108 418
rect 50 130 62 406
rect 96 130 108 406
rect 50 118 108 130
rect -108 -130 -50 -118
rect -108 -406 -96 -130
rect -62 -406 -50 -130
rect -108 -418 -50 -406
rect 50 -130 108 -118
rect 50 -406 62 -130
rect 96 -406 108 -130
rect 50 -418 108 -406
<< pdiffc >>
rect -96 130 -62 406
rect 62 130 96 406
rect -96 -406 -62 -130
rect 62 -406 96 -130
<< nsubdiff >>
rect -210 567 -114 601
rect 114 567 210 601
rect -210 505 -176 567
rect 176 505 210 567
rect -210 -567 -176 -505
rect 176 -567 210 -505
rect -210 -601 -114 -567
rect 114 -601 210 -567
<< nsubdiffcont >>
rect -114 567 114 601
rect -210 -505 -176 505
rect 176 -505 210 505
rect -114 -601 114 -567
<< poly >>
rect -50 499 50 515
rect -50 465 -34 499
rect 34 465 50 499
rect -50 418 50 465
rect -50 71 50 118
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -118 50 -71
rect -50 -465 50 -418
rect -50 -499 -34 -465
rect 34 -499 50 -465
rect -50 -515 50 -499
<< polycont >>
rect -34 465 34 499
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -499 34 -465
<< locali >>
rect -210 567 -114 601
rect 114 567 210 601
rect -210 505 -176 567
rect 176 505 210 567
rect -50 465 -34 499
rect 34 465 50 499
rect -96 406 -62 422
rect -96 114 -62 130
rect 62 406 96 422
rect 62 114 96 130
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -130 -62 -114
rect -96 -422 -62 -406
rect 62 -130 96 -114
rect 62 -422 96 -406
rect -50 -499 -34 -465
rect 34 -499 50 -465
rect -210 -567 -176 -505
rect 176 -567 210 -505
rect -210 -601 -114 -567
rect 114 -601 210 -567
<< viali >>
rect -34 465 34 499
rect -96 130 -62 406
rect 62 130 96 406
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -406 -62 -130
rect 62 -406 96 -130
rect -34 -499 34 -465
<< metal1 >>
rect -46 499 46 505
rect -46 465 -34 499
rect 34 465 46 499
rect -46 459 46 465
rect -102 406 -56 418
rect -102 130 -96 406
rect -62 130 -56 406
rect -102 118 -56 130
rect 56 406 102 418
rect 56 130 62 406
rect 96 130 102 406
rect 56 118 102 130
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -130 -56 -118
rect -102 -406 -96 -130
rect -62 -406 -56 -130
rect -102 -418 -56 -406
rect 56 -130 102 -118
rect 56 -406 62 -130
rect 96 -406 102 -130
rect 56 -418 102 -406
rect -46 -465 46 -459
rect -46 -499 -34 -465
rect 34 -499 46 -465
rect -46 -505 46 -499
<< properties >>
string FIXED_BBOX -193 -584 193 584
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.5 l 0.5 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
