magic
tech sky130A
magscale 1 2
timestamp 1730459124
<< metal3 >>
rect -386 1292 386 1320
rect -386 868 302 1292
rect 366 868 386 1292
rect -386 840 386 868
rect -386 572 386 600
rect -386 148 302 572
rect 366 148 386 572
rect -386 120 386 148
rect -386 -148 386 -120
rect -386 -572 302 -148
rect 366 -572 386 -148
rect -386 -600 386 -572
rect -386 -868 386 -840
rect -386 -1292 302 -868
rect 366 -1292 386 -868
rect -386 -1320 386 -1292
<< via3 >>
rect 302 868 366 1292
rect 302 148 366 572
rect 302 -572 366 -148
rect 302 -1292 366 -868
<< mimcap >>
rect -346 1240 54 1280
rect -346 920 -306 1240
rect 14 920 54 1240
rect -346 880 54 920
rect -346 520 54 560
rect -346 200 -306 520
rect 14 200 54 520
rect -346 160 54 200
rect -346 -200 54 -160
rect -346 -520 -306 -200
rect 14 -520 54 -200
rect -346 -560 54 -520
rect -346 -920 54 -880
rect -346 -1240 -306 -920
rect 14 -1240 54 -920
rect -346 -1280 54 -1240
<< mimcapcontact >>
rect -306 920 14 1240
rect -306 200 14 520
rect -306 -520 14 -200
rect -306 -1240 14 -920
<< metal4 >>
rect -198 1241 -94 1440
rect 282 1292 386 1440
rect -307 1240 15 1241
rect -307 920 -306 1240
rect 14 920 15 1240
rect -307 919 15 920
rect -198 521 -94 919
rect 282 868 302 1292
rect 366 868 386 1292
rect 282 572 386 868
rect -307 520 15 521
rect -307 200 -306 520
rect 14 200 15 520
rect -307 199 15 200
rect -198 -199 -94 199
rect 282 148 302 572
rect 366 148 386 572
rect 282 -148 386 148
rect -307 -200 15 -199
rect -307 -520 -306 -200
rect 14 -520 15 -200
rect -307 -521 15 -520
rect -198 -919 -94 -521
rect 282 -572 302 -148
rect 366 -572 386 -148
rect 282 -868 386 -572
rect -307 -920 15 -919
rect -307 -1240 -306 -920
rect 14 -1240 15 -920
rect -307 -1241 15 -1240
rect -198 -1440 -94 -1241
rect 282 -1292 302 -868
rect 366 -1292 386 -868
rect 282 -1440 386 -1292
<< properties >>
string FIXED_BBOX -386 840 94 1320
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
