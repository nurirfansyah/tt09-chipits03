magic
tech sky130A
magscale 1 2
timestamp 1731265361
<< nwell >>
rect -1696 -819 1696 819
<< pmoslvt >>
rect -1500 -600 1500 600
<< pdiff >>
rect -1558 561 -1500 600
rect -1558 527 -1546 561
rect -1512 527 -1500 561
rect -1558 493 -1500 527
rect -1558 459 -1546 493
rect -1512 459 -1500 493
rect -1558 425 -1500 459
rect -1558 391 -1546 425
rect -1512 391 -1500 425
rect -1558 357 -1500 391
rect -1558 323 -1546 357
rect -1512 323 -1500 357
rect -1558 289 -1500 323
rect -1558 255 -1546 289
rect -1512 255 -1500 289
rect -1558 221 -1500 255
rect -1558 187 -1546 221
rect -1512 187 -1500 221
rect -1558 153 -1500 187
rect -1558 119 -1546 153
rect -1512 119 -1500 153
rect -1558 85 -1500 119
rect -1558 51 -1546 85
rect -1512 51 -1500 85
rect -1558 17 -1500 51
rect -1558 -17 -1546 17
rect -1512 -17 -1500 17
rect -1558 -51 -1500 -17
rect -1558 -85 -1546 -51
rect -1512 -85 -1500 -51
rect -1558 -119 -1500 -85
rect -1558 -153 -1546 -119
rect -1512 -153 -1500 -119
rect -1558 -187 -1500 -153
rect -1558 -221 -1546 -187
rect -1512 -221 -1500 -187
rect -1558 -255 -1500 -221
rect -1558 -289 -1546 -255
rect -1512 -289 -1500 -255
rect -1558 -323 -1500 -289
rect -1558 -357 -1546 -323
rect -1512 -357 -1500 -323
rect -1558 -391 -1500 -357
rect -1558 -425 -1546 -391
rect -1512 -425 -1500 -391
rect -1558 -459 -1500 -425
rect -1558 -493 -1546 -459
rect -1512 -493 -1500 -459
rect -1558 -527 -1500 -493
rect -1558 -561 -1546 -527
rect -1512 -561 -1500 -527
rect -1558 -600 -1500 -561
rect 1500 561 1558 600
rect 1500 527 1512 561
rect 1546 527 1558 561
rect 1500 493 1558 527
rect 1500 459 1512 493
rect 1546 459 1558 493
rect 1500 425 1558 459
rect 1500 391 1512 425
rect 1546 391 1558 425
rect 1500 357 1558 391
rect 1500 323 1512 357
rect 1546 323 1558 357
rect 1500 289 1558 323
rect 1500 255 1512 289
rect 1546 255 1558 289
rect 1500 221 1558 255
rect 1500 187 1512 221
rect 1546 187 1558 221
rect 1500 153 1558 187
rect 1500 119 1512 153
rect 1546 119 1558 153
rect 1500 85 1558 119
rect 1500 51 1512 85
rect 1546 51 1558 85
rect 1500 17 1558 51
rect 1500 -17 1512 17
rect 1546 -17 1558 17
rect 1500 -51 1558 -17
rect 1500 -85 1512 -51
rect 1546 -85 1558 -51
rect 1500 -119 1558 -85
rect 1500 -153 1512 -119
rect 1546 -153 1558 -119
rect 1500 -187 1558 -153
rect 1500 -221 1512 -187
rect 1546 -221 1558 -187
rect 1500 -255 1558 -221
rect 1500 -289 1512 -255
rect 1546 -289 1558 -255
rect 1500 -323 1558 -289
rect 1500 -357 1512 -323
rect 1546 -357 1558 -323
rect 1500 -391 1558 -357
rect 1500 -425 1512 -391
rect 1546 -425 1558 -391
rect 1500 -459 1558 -425
rect 1500 -493 1512 -459
rect 1546 -493 1558 -459
rect 1500 -527 1558 -493
rect 1500 -561 1512 -527
rect 1546 -561 1558 -527
rect 1500 -600 1558 -561
<< pdiffc >>
rect -1546 527 -1512 561
rect -1546 459 -1512 493
rect -1546 391 -1512 425
rect -1546 323 -1512 357
rect -1546 255 -1512 289
rect -1546 187 -1512 221
rect -1546 119 -1512 153
rect -1546 51 -1512 85
rect -1546 -17 -1512 17
rect -1546 -85 -1512 -51
rect -1546 -153 -1512 -119
rect -1546 -221 -1512 -187
rect -1546 -289 -1512 -255
rect -1546 -357 -1512 -323
rect -1546 -425 -1512 -391
rect -1546 -493 -1512 -459
rect -1546 -561 -1512 -527
rect 1512 527 1546 561
rect 1512 459 1546 493
rect 1512 391 1546 425
rect 1512 323 1546 357
rect 1512 255 1546 289
rect 1512 187 1546 221
rect 1512 119 1546 153
rect 1512 51 1546 85
rect 1512 -17 1546 17
rect 1512 -85 1546 -51
rect 1512 -153 1546 -119
rect 1512 -221 1546 -187
rect 1512 -289 1546 -255
rect 1512 -357 1546 -323
rect 1512 -425 1546 -391
rect 1512 -493 1546 -459
rect 1512 -561 1546 -527
<< nsubdiff >>
rect -1660 749 -1547 783
rect -1513 749 -1479 783
rect -1445 749 -1411 783
rect -1377 749 -1343 783
rect -1309 749 -1275 783
rect -1241 749 -1207 783
rect -1173 749 -1139 783
rect -1105 749 -1071 783
rect -1037 749 -1003 783
rect -969 749 -935 783
rect -901 749 -867 783
rect -833 749 -799 783
rect -765 749 -731 783
rect -697 749 -663 783
rect -629 749 -595 783
rect -561 749 -527 783
rect -493 749 -459 783
rect -425 749 -391 783
rect -357 749 -323 783
rect -289 749 -255 783
rect -221 749 -187 783
rect -153 749 -119 783
rect -85 749 -51 783
rect -17 749 17 783
rect 51 749 85 783
rect 119 749 153 783
rect 187 749 221 783
rect 255 749 289 783
rect 323 749 357 783
rect 391 749 425 783
rect 459 749 493 783
rect 527 749 561 783
rect 595 749 629 783
rect 663 749 697 783
rect 731 749 765 783
rect 799 749 833 783
rect 867 749 901 783
rect 935 749 969 783
rect 1003 749 1037 783
rect 1071 749 1105 783
rect 1139 749 1173 783
rect 1207 749 1241 783
rect 1275 749 1309 783
rect 1343 749 1377 783
rect 1411 749 1445 783
rect 1479 749 1513 783
rect 1547 749 1660 783
rect -1660 663 -1626 749
rect -1660 595 -1626 629
rect 1626 663 1660 749
rect -1660 527 -1626 561
rect -1660 459 -1626 493
rect -1660 391 -1626 425
rect -1660 323 -1626 357
rect -1660 255 -1626 289
rect -1660 187 -1626 221
rect -1660 119 -1626 153
rect -1660 51 -1626 85
rect -1660 -17 -1626 17
rect -1660 -85 -1626 -51
rect -1660 -153 -1626 -119
rect -1660 -221 -1626 -187
rect -1660 -289 -1626 -255
rect -1660 -357 -1626 -323
rect -1660 -425 -1626 -391
rect -1660 -493 -1626 -459
rect -1660 -561 -1626 -527
rect -1660 -629 -1626 -595
rect 1626 595 1660 629
rect 1626 527 1660 561
rect 1626 459 1660 493
rect 1626 391 1660 425
rect 1626 323 1660 357
rect 1626 255 1660 289
rect 1626 187 1660 221
rect 1626 119 1660 153
rect 1626 51 1660 85
rect 1626 -17 1660 17
rect 1626 -85 1660 -51
rect 1626 -153 1660 -119
rect 1626 -221 1660 -187
rect 1626 -289 1660 -255
rect 1626 -357 1660 -323
rect 1626 -425 1660 -391
rect 1626 -493 1660 -459
rect 1626 -561 1660 -527
rect -1660 -749 -1626 -663
rect 1626 -629 1660 -595
rect 1626 -749 1660 -663
rect -1660 -783 -1547 -749
rect -1513 -783 -1479 -749
rect -1445 -783 -1411 -749
rect -1377 -783 -1343 -749
rect -1309 -783 -1275 -749
rect -1241 -783 -1207 -749
rect -1173 -783 -1139 -749
rect -1105 -783 -1071 -749
rect -1037 -783 -1003 -749
rect -969 -783 -935 -749
rect -901 -783 -867 -749
rect -833 -783 -799 -749
rect -765 -783 -731 -749
rect -697 -783 -663 -749
rect -629 -783 -595 -749
rect -561 -783 -527 -749
rect -493 -783 -459 -749
rect -425 -783 -391 -749
rect -357 -783 -323 -749
rect -289 -783 -255 -749
rect -221 -783 -187 -749
rect -153 -783 -119 -749
rect -85 -783 -51 -749
rect -17 -783 17 -749
rect 51 -783 85 -749
rect 119 -783 153 -749
rect 187 -783 221 -749
rect 255 -783 289 -749
rect 323 -783 357 -749
rect 391 -783 425 -749
rect 459 -783 493 -749
rect 527 -783 561 -749
rect 595 -783 629 -749
rect 663 -783 697 -749
rect 731 -783 765 -749
rect 799 -783 833 -749
rect 867 -783 901 -749
rect 935 -783 969 -749
rect 1003 -783 1037 -749
rect 1071 -783 1105 -749
rect 1139 -783 1173 -749
rect 1207 -783 1241 -749
rect 1275 -783 1309 -749
rect 1343 -783 1377 -749
rect 1411 -783 1445 -749
rect 1479 -783 1513 -749
rect 1547 -783 1660 -749
<< nsubdiffcont >>
rect -1547 749 -1513 783
rect -1479 749 -1445 783
rect -1411 749 -1377 783
rect -1343 749 -1309 783
rect -1275 749 -1241 783
rect -1207 749 -1173 783
rect -1139 749 -1105 783
rect -1071 749 -1037 783
rect -1003 749 -969 783
rect -935 749 -901 783
rect -867 749 -833 783
rect -799 749 -765 783
rect -731 749 -697 783
rect -663 749 -629 783
rect -595 749 -561 783
rect -527 749 -493 783
rect -459 749 -425 783
rect -391 749 -357 783
rect -323 749 -289 783
rect -255 749 -221 783
rect -187 749 -153 783
rect -119 749 -85 783
rect -51 749 -17 783
rect 17 749 51 783
rect 85 749 119 783
rect 153 749 187 783
rect 221 749 255 783
rect 289 749 323 783
rect 357 749 391 783
rect 425 749 459 783
rect 493 749 527 783
rect 561 749 595 783
rect 629 749 663 783
rect 697 749 731 783
rect 765 749 799 783
rect 833 749 867 783
rect 901 749 935 783
rect 969 749 1003 783
rect 1037 749 1071 783
rect 1105 749 1139 783
rect 1173 749 1207 783
rect 1241 749 1275 783
rect 1309 749 1343 783
rect 1377 749 1411 783
rect 1445 749 1479 783
rect 1513 749 1547 783
rect -1660 629 -1626 663
rect 1626 629 1660 663
rect -1660 561 -1626 595
rect -1660 493 -1626 527
rect -1660 425 -1626 459
rect -1660 357 -1626 391
rect -1660 289 -1626 323
rect -1660 221 -1626 255
rect -1660 153 -1626 187
rect -1660 85 -1626 119
rect -1660 17 -1626 51
rect -1660 -51 -1626 -17
rect -1660 -119 -1626 -85
rect -1660 -187 -1626 -153
rect -1660 -255 -1626 -221
rect -1660 -323 -1626 -289
rect -1660 -391 -1626 -357
rect -1660 -459 -1626 -425
rect -1660 -527 -1626 -493
rect -1660 -595 -1626 -561
rect 1626 561 1660 595
rect 1626 493 1660 527
rect 1626 425 1660 459
rect 1626 357 1660 391
rect 1626 289 1660 323
rect 1626 221 1660 255
rect 1626 153 1660 187
rect 1626 85 1660 119
rect 1626 17 1660 51
rect 1626 -51 1660 -17
rect 1626 -119 1660 -85
rect 1626 -187 1660 -153
rect 1626 -255 1660 -221
rect 1626 -323 1660 -289
rect 1626 -391 1660 -357
rect 1626 -459 1660 -425
rect 1626 -527 1660 -493
rect 1626 -595 1660 -561
rect -1660 -663 -1626 -629
rect 1626 -663 1660 -629
rect -1547 -783 -1513 -749
rect -1479 -783 -1445 -749
rect -1411 -783 -1377 -749
rect -1343 -783 -1309 -749
rect -1275 -783 -1241 -749
rect -1207 -783 -1173 -749
rect -1139 -783 -1105 -749
rect -1071 -783 -1037 -749
rect -1003 -783 -969 -749
rect -935 -783 -901 -749
rect -867 -783 -833 -749
rect -799 -783 -765 -749
rect -731 -783 -697 -749
rect -663 -783 -629 -749
rect -595 -783 -561 -749
rect -527 -783 -493 -749
rect -459 -783 -425 -749
rect -391 -783 -357 -749
rect -323 -783 -289 -749
rect -255 -783 -221 -749
rect -187 -783 -153 -749
rect -119 -783 -85 -749
rect -51 -783 -17 -749
rect 17 -783 51 -749
rect 85 -783 119 -749
rect 153 -783 187 -749
rect 221 -783 255 -749
rect 289 -783 323 -749
rect 357 -783 391 -749
rect 425 -783 459 -749
rect 493 -783 527 -749
rect 561 -783 595 -749
rect 629 -783 663 -749
rect 697 -783 731 -749
rect 765 -783 799 -749
rect 833 -783 867 -749
rect 901 -783 935 -749
rect 969 -783 1003 -749
rect 1037 -783 1071 -749
rect 1105 -783 1139 -749
rect 1173 -783 1207 -749
rect 1241 -783 1275 -749
rect 1309 -783 1343 -749
rect 1377 -783 1411 -749
rect 1445 -783 1479 -749
rect 1513 -783 1547 -749
<< poly >>
rect -1500 681 1500 697
rect -1500 647 -1479 681
rect -1445 647 -1411 681
rect -1377 647 -1343 681
rect -1309 647 -1275 681
rect -1241 647 -1207 681
rect -1173 647 -1139 681
rect -1105 647 -1071 681
rect -1037 647 -1003 681
rect -969 647 -935 681
rect -901 647 -867 681
rect -833 647 -799 681
rect -765 647 -731 681
rect -697 647 -663 681
rect -629 647 -595 681
rect -561 647 -527 681
rect -493 647 -459 681
rect -425 647 -391 681
rect -357 647 -323 681
rect -289 647 -255 681
rect -221 647 -187 681
rect -153 647 -119 681
rect -85 647 -51 681
rect -17 647 17 681
rect 51 647 85 681
rect 119 647 153 681
rect 187 647 221 681
rect 255 647 289 681
rect 323 647 357 681
rect 391 647 425 681
rect 459 647 493 681
rect 527 647 561 681
rect 595 647 629 681
rect 663 647 697 681
rect 731 647 765 681
rect 799 647 833 681
rect 867 647 901 681
rect 935 647 969 681
rect 1003 647 1037 681
rect 1071 647 1105 681
rect 1139 647 1173 681
rect 1207 647 1241 681
rect 1275 647 1309 681
rect 1343 647 1377 681
rect 1411 647 1445 681
rect 1479 647 1500 681
rect -1500 600 1500 647
rect -1500 -647 1500 -600
rect -1500 -681 -1479 -647
rect -1445 -681 -1411 -647
rect -1377 -681 -1343 -647
rect -1309 -681 -1275 -647
rect -1241 -681 -1207 -647
rect -1173 -681 -1139 -647
rect -1105 -681 -1071 -647
rect -1037 -681 -1003 -647
rect -969 -681 -935 -647
rect -901 -681 -867 -647
rect -833 -681 -799 -647
rect -765 -681 -731 -647
rect -697 -681 -663 -647
rect -629 -681 -595 -647
rect -561 -681 -527 -647
rect -493 -681 -459 -647
rect -425 -681 -391 -647
rect -357 -681 -323 -647
rect -289 -681 -255 -647
rect -221 -681 -187 -647
rect -153 -681 -119 -647
rect -85 -681 -51 -647
rect -17 -681 17 -647
rect 51 -681 85 -647
rect 119 -681 153 -647
rect 187 -681 221 -647
rect 255 -681 289 -647
rect 323 -681 357 -647
rect 391 -681 425 -647
rect 459 -681 493 -647
rect 527 -681 561 -647
rect 595 -681 629 -647
rect 663 -681 697 -647
rect 731 -681 765 -647
rect 799 -681 833 -647
rect 867 -681 901 -647
rect 935 -681 969 -647
rect 1003 -681 1037 -647
rect 1071 -681 1105 -647
rect 1139 -681 1173 -647
rect 1207 -681 1241 -647
rect 1275 -681 1309 -647
rect 1343 -681 1377 -647
rect 1411 -681 1445 -647
rect 1479 -681 1500 -647
rect -1500 -697 1500 -681
<< polycont >>
rect -1479 647 -1445 681
rect -1411 647 -1377 681
rect -1343 647 -1309 681
rect -1275 647 -1241 681
rect -1207 647 -1173 681
rect -1139 647 -1105 681
rect -1071 647 -1037 681
rect -1003 647 -969 681
rect -935 647 -901 681
rect -867 647 -833 681
rect -799 647 -765 681
rect -731 647 -697 681
rect -663 647 -629 681
rect -595 647 -561 681
rect -527 647 -493 681
rect -459 647 -425 681
rect -391 647 -357 681
rect -323 647 -289 681
rect -255 647 -221 681
rect -187 647 -153 681
rect -119 647 -85 681
rect -51 647 -17 681
rect 17 647 51 681
rect 85 647 119 681
rect 153 647 187 681
rect 221 647 255 681
rect 289 647 323 681
rect 357 647 391 681
rect 425 647 459 681
rect 493 647 527 681
rect 561 647 595 681
rect 629 647 663 681
rect 697 647 731 681
rect 765 647 799 681
rect 833 647 867 681
rect 901 647 935 681
rect 969 647 1003 681
rect 1037 647 1071 681
rect 1105 647 1139 681
rect 1173 647 1207 681
rect 1241 647 1275 681
rect 1309 647 1343 681
rect 1377 647 1411 681
rect 1445 647 1479 681
rect -1479 -681 -1445 -647
rect -1411 -681 -1377 -647
rect -1343 -681 -1309 -647
rect -1275 -681 -1241 -647
rect -1207 -681 -1173 -647
rect -1139 -681 -1105 -647
rect -1071 -681 -1037 -647
rect -1003 -681 -969 -647
rect -935 -681 -901 -647
rect -867 -681 -833 -647
rect -799 -681 -765 -647
rect -731 -681 -697 -647
rect -663 -681 -629 -647
rect -595 -681 -561 -647
rect -527 -681 -493 -647
rect -459 -681 -425 -647
rect -391 -681 -357 -647
rect -323 -681 -289 -647
rect -255 -681 -221 -647
rect -187 -681 -153 -647
rect -119 -681 -85 -647
rect -51 -681 -17 -647
rect 17 -681 51 -647
rect 85 -681 119 -647
rect 153 -681 187 -647
rect 221 -681 255 -647
rect 289 -681 323 -647
rect 357 -681 391 -647
rect 425 -681 459 -647
rect 493 -681 527 -647
rect 561 -681 595 -647
rect 629 -681 663 -647
rect 697 -681 731 -647
rect 765 -681 799 -647
rect 833 -681 867 -647
rect 901 -681 935 -647
rect 969 -681 1003 -647
rect 1037 -681 1071 -647
rect 1105 -681 1139 -647
rect 1173 -681 1207 -647
rect 1241 -681 1275 -647
rect 1309 -681 1343 -647
rect 1377 -681 1411 -647
rect 1445 -681 1479 -647
<< locali >>
rect -1660 749 -1547 783
rect -1513 749 -1479 783
rect -1445 749 -1411 783
rect -1377 749 -1343 783
rect -1309 749 -1275 783
rect -1241 749 -1207 783
rect -1173 749 -1139 783
rect -1105 749 -1071 783
rect -1037 749 -1003 783
rect -969 749 -935 783
rect -901 749 -867 783
rect -833 749 -799 783
rect -765 749 -731 783
rect -697 749 -663 783
rect -629 749 -595 783
rect -561 749 -527 783
rect -493 749 -459 783
rect -425 749 -391 783
rect -357 749 -323 783
rect -289 749 -255 783
rect -221 749 -187 783
rect -153 749 -119 783
rect -85 749 -51 783
rect -17 749 17 783
rect 51 749 85 783
rect 119 749 153 783
rect 187 749 221 783
rect 255 749 289 783
rect 323 749 357 783
rect 391 749 425 783
rect 459 749 493 783
rect 527 749 561 783
rect 595 749 629 783
rect 663 749 697 783
rect 731 749 765 783
rect 799 749 833 783
rect 867 749 901 783
rect 935 749 969 783
rect 1003 749 1037 783
rect 1071 749 1105 783
rect 1139 749 1173 783
rect 1207 749 1241 783
rect 1275 749 1309 783
rect 1343 749 1377 783
rect 1411 749 1445 783
rect 1479 749 1513 783
rect 1547 749 1660 783
rect -1660 663 -1626 749
rect -1500 647 -1479 681
rect -1423 647 -1411 681
rect -1351 647 -1343 681
rect -1279 647 -1275 681
rect -1173 647 -1169 681
rect -1105 647 -1097 681
rect -1037 647 -1025 681
rect -969 647 -953 681
rect -901 647 -881 681
rect -833 647 -809 681
rect -765 647 -737 681
rect -697 647 -665 681
rect -629 647 -595 681
rect -559 647 -527 681
rect -487 647 -459 681
rect -415 647 -391 681
rect -343 647 -323 681
rect -271 647 -255 681
rect -199 647 -187 681
rect -127 647 -119 681
rect -55 647 -51 681
rect 51 647 55 681
rect 119 647 127 681
rect 187 647 199 681
rect 255 647 271 681
rect 323 647 343 681
rect 391 647 415 681
rect 459 647 487 681
rect 527 647 559 681
rect 595 647 629 681
rect 665 647 697 681
rect 737 647 765 681
rect 809 647 833 681
rect 881 647 901 681
rect 953 647 969 681
rect 1025 647 1037 681
rect 1097 647 1105 681
rect 1169 647 1173 681
rect 1275 647 1279 681
rect 1343 647 1351 681
rect 1411 647 1423 681
rect 1479 647 1500 681
rect 1626 663 1660 749
rect -1660 595 -1626 629
rect -1660 527 -1626 561
rect -1660 459 -1626 493
rect -1660 391 -1626 425
rect -1660 323 -1626 357
rect -1660 255 -1626 289
rect -1660 187 -1626 221
rect -1660 119 -1626 153
rect -1660 51 -1626 85
rect -1660 -17 -1626 17
rect -1660 -85 -1626 -51
rect -1660 -153 -1626 -119
rect -1660 -221 -1626 -187
rect -1660 -289 -1626 -255
rect -1660 -357 -1626 -323
rect -1660 -425 -1626 -391
rect -1660 -493 -1626 -459
rect -1660 -561 -1626 -527
rect -1660 -629 -1626 -595
rect -1546 561 -1512 604
rect -1546 493 -1512 523
rect -1546 425 -1512 451
rect -1546 357 -1512 379
rect -1546 289 -1512 307
rect -1546 221 -1512 235
rect -1546 153 -1512 163
rect -1546 85 -1512 91
rect -1546 17 -1512 19
rect -1546 -19 -1512 -17
rect -1546 -91 -1512 -85
rect -1546 -163 -1512 -153
rect -1546 -235 -1512 -221
rect -1546 -307 -1512 -289
rect -1546 -379 -1512 -357
rect -1546 -451 -1512 -425
rect -1546 -523 -1512 -493
rect -1546 -604 -1512 -561
rect 1512 561 1546 604
rect 1512 493 1546 523
rect 1512 425 1546 451
rect 1512 357 1546 379
rect 1512 289 1546 307
rect 1512 221 1546 235
rect 1512 153 1546 163
rect 1512 85 1546 91
rect 1512 17 1546 19
rect 1512 -19 1546 -17
rect 1512 -91 1546 -85
rect 1512 -163 1546 -153
rect 1512 -235 1546 -221
rect 1512 -307 1546 -289
rect 1512 -379 1546 -357
rect 1512 -451 1546 -425
rect 1512 -523 1546 -493
rect 1512 -604 1546 -561
rect 1626 595 1660 629
rect 1626 527 1660 561
rect 1626 459 1660 493
rect 1626 391 1660 425
rect 1626 323 1660 357
rect 1626 255 1660 289
rect 1626 187 1660 221
rect 1626 119 1660 153
rect 1626 51 1660 85
rect 1626 -17 1660 17
rect 1626 -85 1660 -51
rect 1626 -153 1660 -119
rect 1626 -221 1660 -187
rect 1626 -289 1660 -255
rect 1626 -357 1660 -323
rect 1626 -425 1660 -391
rect 1626 -493 1660 -459
rect 1626 -561 1660 -527
rect 1626 -629 1660 -595
rect -1660 -749 -1626 -663
rect -1500 -681 -1479 -647
rect -1423 -681 -1411 -647
rect -1351 -681 -1343 -647
rect -1279 -681 -1275 -647
rect -1173 -681 -1169 -647
rect -1105 -681 -1097 -647
rect -1037 -681 -1025 -647
rect -969 -681 -953 -647
rect -901 -681 -881 -647
rect -833 -681 -809 -647
rect -765 -681 -737 -647
rect -697 -681 -665 -647
rect -629 -681 -595 -647
rect -559 -681 -527 -647
rect -487 -681 -459 -647
rect -415 -681 -391 -647
rect -343 -681 -323 -647
rect -271 -681 -255 -647
rect -199 -681 -187 -647
rect -127 -681 -119 -647
rect -55 -681 -51 -647
rect 51 -681 55 -647
rect 119 -681 127 -647
rect 187 -681 199 -647
rect 255 -681 271 -647
rect 323 -681 343 -647
rect 391 -681 415 -647
rect 459 -681 487 -647
rect 527 -681 559 -647
rect 595 -681 629 -647
rect 665 -681 697 -647
rect 737 -681 765 -647
rect 809 -681 833 -647
rect 881 -681 901 -647
rect 953 -681 969 -647
rect 1025 -681 1037 -647
rect 1097 -681 1105 -647
rect 1169 -681 1173 -647
rect 1275 -681 1279 -647
rect 1343 -681 1351 -647
rect 1411 -681 1423 -647
rect 1479 -681 1500 -647
rect 1626 -749 1660 -663
rect -1660 -783 -1547 -749
rect -1513 -783 -1479 -749
rect -1445 -783 -1411 -749
rect -1377 -783 -1343 -749
rect -1309 -783 -1275 -749
rect -1241 -783 -1207 -749
rect -1173 -783 -1139 -749
rect -1105 -783 -1071 -749
rect -1037 -783 -1003 -749
rect -969 -783 -935 -749
rect -901 -783 -867 -749
rect -833 -783 -799 -749
rect -765 -783 -731 -749
rect -697 -783 -663 -749
rect -629 -783 -595 -749
rect -561 -783 -527 -749
rect -493 -783 -459 -749
rect -425 -783 -391 -749
rect -357 -783 -323 -749
rect -289 -783 -255 -749
rect -221 -783 -187 -749
rect -153 -783 -119 -749
rect -85 -783 -51 -749
rect -17 -783 17 -749
rect 51 -783 85 -749
rect 119 -783 153 -749
rect 187 -783 221 -749
rect 255 -783 289 -749
rect 323 -783 357 -749
rect 391 -783 425 -749
rect 459 -783 493 -749
rect 527 -783 561 -749
rect 595 -783 629 -749
rect 663 -783 697 -749
rect 731 -783 765 -749
rect 799 -783 833 -749
rect 867 -783 901 -749
rect 935 -783 969 -749
rect 1003 -783 1037 -749
rect 1071 -783 1105 -749
rect 1139 -783 1173 -749
rect 1207 -783 1241 -749
rect 1275 -783 1309 -749
rect 1343 -783 1377 -749
rect 1411 -783 1445 -749
rect 1479 -783 1513 -749
rect 1547 -783 1660 -749
<< viali >>
rect -1457 647 -1445 681
rect -1445 647 -1423 681
rect -1385 647 -1377 681
rect -1377 647 -1351 681
rect -1313 647 -1309 681
rect -1309 647 -1279 681
rect -1241 647 -1207 681
rect -1169 647 -1139 681
rect -1139 647 -1135 681
rect -1097 647 -1071 681
rect -1071 647 -1063 681
rect -1025 647 -1003 681
rect -1003 647 -991 681
rect -953 647 -935 681
rect -935 647 -919 681
rect -881 647 -867 681
rect -867 647 -847 681
rect -809 647 -799 681
rect -799 647 -775 681
rect -737 647 -731 681
rect -731 647 -703 681
rect -665 647 -663 681
rect -663 647 -631 681
rect -593 647 -561 681
rect -561 647 -559 681
rect -521 647 -493 681
rect -493 647 -487 681
rect -449 647 -425 681
rect -425 647 -415 681
rect -377 647 -357 681
rect -357 647 -343 681
rect -305 647 -289 681
rect -289 647 -271 681
rect -233 647 -221 681
rect -221 647 -199 681
rect -161 647 -153 681
rect -153 647 -127 681
rect -89 647 -85 681
rect -85 647 -55 681
rect -17 647 17 681
rect 55 647 85 681
rect 85 647 89 681
rect 127 647 153 681
rect 153 647 161 681
rect 199 647 221 681
rect 221 647 233 681
rect 271 647 289 681
rect 289 647 305 681
rect 343 647 357 681
rect 357 647 377 681
rect 415 647 425 681
rect 425 647 449 681
rect 487 647 493 681
rect 493 647 521 681
rect 559 647 561 681
rect 561 647 593 681
rect 631 647 663 681
rect 663 647 665 681
rect 703 647 731 681
rect 731 647 737 681
rect 775 647 799 681
rect 799 647 809 681
rect 847 647 867 681
rect 867 647 881 681
rect 919 647 935 681
rect 935 647 953 681
rect 991 647 1003 681
rect 1003 647 1025 681
rect 1063 647 1071 681
rect 1071 647 1097 681
rect 1135 647 1139 681
rect 1139 647 1169 681
rect 1207 647 1241 681
rect 1279 647 1309 681
rect 1309 647 1313 681
rect 1351 647 1377 681
rect 1377 647 1385 681
rect 1423 647 1445 681
rect 1445 647 1457 681
rect -1546 527 -1512 557
rect -1546 523 -1512 527
rect -1546 459 -1512 485
rect -1546 451 -1512 459
rect -1546 391 -1512 413
rect -1546 379 -1512 391
rect -1546 323 -1512 341
rect -1546 307 -1512 323
rect -1546 255 -1512 269
rect -1546 235 -1512 255
rect -1546 187 -1512 197
rect -1546 163 -1512 187
rect -1546 119 -1512 125
rect -1546 91 -1512 119
rect -1546 51 -1512 53
rect -1546 19 -1512 51
rect -1546 -51 -1512 -19
rect -1546 -53 -1512 -51
rect -1546 -119 -1512 -91
rect -1546 -125 -1512 -119
rect -1546 -187 -1512 -163
rect -1546 -197 -1512 -187
rect -1546 -255 -1512 -235
rect -1546 -269 -1512 -255
rect -1546 -323 -1512 -307
rect -1546 -341 -1512 -323
rect -1546 -391 -1512 -379
rect -1546 -413 -1512 -391
rect -1546 -459 -1512 -451
rect -1546 -485 -1512 -459
rect -1546 -527 -1512 -523
rect -1546 -557 -1512 -527
rect 1512 527 1546 557
rect 1512 523 1546 527
rect 1512 459 1546 485
rect 1512 451 1546 459
rect 1512 391 1546 413
rect 1512 379 1546 391
rect 1512 323 1546 341
rect 1512 307 1546 323
rect 1512 255 1546 269
rect 1512 235 1546 255
rect 1512 187 1546 197
rect 1512 163 1546 187
rect 1512 119 1546 125
rect 1512 91 1546 119
rect 1512 51 1546 53
rect 1512 19 1546 51
rect 1512 -51 1546 -19
rect 1512 -53 1546 -51
rect 1512 -119 1546 -91
rect 1512 -125 1546 -119
rect 1512 -187 1546 -163
rect 1512 -197 1546 -187
rect 1512 -255 1546 -235
rect 1512 -269 1546 -255
rect 1512 -323 1546 -307
rect 1512 -341 1546 -323
rect 1512 -391 1546 -379
rect 1512 -413 1546 -391
rect 1512 -459 1546 -451
rect 1512 -485 1546 -459
rect 1512 -527 1546 -523
rect 1512 -557 1546 -527
rect -1457 -681 -1445 -647
rect -1445 -681 -1423 -647
rect -1385 -681 -1377 -647
rect -1377 -681 -1351 -647
rect -1313 -681 -1309 -647
rect -1309 -681 -1279 -647
rect -1241 -681 -1207 -647
rect -1169 -681 -1139 -647
rect -1139 -681 -1135 -647
rect -1097 -681 -1071 -647
rect -1071 -681 -1063 -647
rect -1025 -681 -1003 -647
rect -1003 -681 -991 -647
rect -953 -681 -935 -647
rect -935 -681 -919 -647
rect -881 -681 -867 -647
rect -867 -681 -847 -647
rect -809 -681 -799 -647
rect -799 -681 -775 -647
rect -737 -681 -731 -647
rect -731 -681 -703 -647
rect -665 -681 -663 -647
rect -663 -681 -631 -647
rect -593 -681 -561 -647
rect -561 -681 -559 -647
rect -521 -681 -493 -647
rect -493 -681 -487 -647
rect -449 -681 -425 -647
rect -425 -681 -415 -647
rect -377 -681 -357 -647
rect -357 -681 -343 -647
rect -305 -681 -289 -647
rect -289 -681 -271 -647
rect -233 -681 -221 -647
rect -221 -681 -199 -647
rect -161 -681 -153 -647
rect -153 -681 -127 -647
rect -89 -681 -85 -647
rect -85 -681 -55 -647
rect -17 -681 17 -647
rect 55 -681 85 -647
rect 85 -681 89 -647
rect 127 -681 153 -647
rect 153 -681 161 -647
rect 199 -681 221 -647
rect 221 -681 233 -647
rect 271 -681 289 -647
rect 289 -681 305 -647
rect 343 -681 357 -647
rect 357 -681 377 -647
rect 415 -681 425 -647
rect 425 -681 449 -647
rect 487 -681 493 -647
rect 493 -681 521 -647
rect 559 -681 561 -647
rect 561 -681 593 -647
rect 631 -681 663 -647
rect 663 -681 665 -647
rect 703 -681 731 -647
rect 731 -681 737 -647
rect 775 -681 799 -647
rect 799 -681 809 -647
rect 847 -681 867 -647
rect 867 -681 881 -647
rect 919 -681 935 -647
rect 935 -681 953 -647
rect 991 -681 1003 -647
rect 1003 -681 1025 -647
rect 1063 -681 1071 -647
rect 1071 -681 1097 -647
rect 1135 -681 1139 -647
rect 1139 -681 1169 -647
rect 1207 -681 1241 -647
rect 1279 -681 1309 -647
rect 1309 -681 1313 -647
rect 1351 -681 1377 -647
rect 1377 -681 1385 -647
rect 1423 -681 1445 -647
rect 1445 -681 1457 -647
<< metal1 >>
rect -1496 681 1496 687
rect -1496 647 -1457 681
rect -1423 647 -1385 681
rect -1351 647 -1313 681
rect -1279 647 -1241 681
rect -1207 647 -1169 681
rect -1135 647 -1097 681
rect -1063 647 -1025 681
rect -991 647 -953 681
rect -919 647 -881 681
rect -847 647 -809 681
rect -775 647 -737 681
rect -703 647 -665 681
rect -631 647 -593 681
rect -559 647 -521 681
rect -487 647 -449 681
rect -415 647 -377 681
rect -343 647 -305 681
rect -271 647 -233 681
rect -199 647 -161 681
rect -127 647 -89 681
rect -55 647 -17 681
rect 17 647 55 681
rect 89 647 127 681
rect 161 647 199 681
rect 233 647 271 681
rect 305 647 343 681
rect 377 647 415 681
rect 449 647 487 681
rect 521 647 559 681
rect 593 647 631 681
rect 665 647 703 681
rect 737 647 775 681
rect 809 647 847 681
rect 881 647 919 681
rect 953 647 991 681
rect 1025 647 1063 681
rect 1097 647 1135 681
rect 1169 647 1207 681
rect 1241 647 1279 681
rect 1313 647 1351 681
rect 1385 647 1423 681
rect 1457 647 1496 681
rect -1496 641 1496 647
rect -1552 557 -1506 600
rect -1552 523 -1546 557
rect -1512 523 -1506 557
rect -1552 485 -1506 523
rect -1552 451 -1546 485
rect -1512 451 -1506 485
rect -1552 413 -1506 451
rect -1552 379 -1546 413
rect -1512 379 -1506 413
rect -1552 341 -1506 379
rect -1552 307 -1546 341
rect -1512 307 -1506 341
rect -1552 269 -1506 307
rect -1552 235 -1546 269
rect -1512 235 -1506 269
rect -1552 197 -1506 235
rect -1552 163 -1546 197
rect -1512 163 -1506 197
rect -1552 125 -1506 163
rect -1552 91 -1546 125
rect -1512 91 -1506 125
rect -1552 53 -1506 91
rect -1552 19 -1546 53
rect -1512 19 -1506 53
rect -1552 -19 -1506 19
rect -1552 -53 -1546 -19
rect -1512 -53 -1506 -19
rect -1552 -91 -1506 -53
rect -1552 -125 -1546 -91
rect -1512 -125 -1506 -91
rect -1552 -163 -1506 -125
rect -1552 -197 -1546 -163
rect -1512 -197 -1506 -163
rect -1552 -235 -1506 -197
rect -1552 -269 -1546 -235
rect -1512 -269 -1506 -235
rect -1552 -307 -1506 -269
rect -1552 -341 -1546 -307
rect -1512 -341 -1506 -307
rect -1552 -379 -1506 -341
rect -1552 -413 -1546 -379
rect -1512 -413 -1506 -379
rect -1552 -451 -1506 -413
rect -1552 -485 -1546 -451
rect -1512 -485 -1506 -451
rect -1552 -523 -1506 -485
rect -1552 -557 -1546 -523
rect -1512 -557 -1506 -523
rect -1552 -600 -1506 -557
rect 1506 557 1552 600
rect 1506 523 1512 557
rect 1546 523 1552 557
rect 1506 485 1552 523
rect 1506 451 1512 485
rect 1546 451 1552 485
rect 1506 413 1552 451
rect 1506 379 1512 413
rect 1546 379 1552 413
rect 1506 341 1552 379
rect 1506 307 1512 341
rect 1546 307 1552 341
rect 1506 269 1552 307
rect 1506 235 1512 269
rect 1546 235 1552 269
rect 1506 197 1552 235
rect 1506 163 1512 197
rect 1546 163 1552 197
rect 1506 125 1552 163
rect 1506 91 1512 125
rect 1546 91 1552 125
rect 1506 53 1552 91
rect 1506 19 1512 53
rect 1546 19 1552 53
rect 1506 -19 1552 19
rect 1506 -53 1512 -19
rect 1546 -53 1552 -19
rect 1506 -91 1552 -53
rect 1506 -125 1512 -91
rect 1546 -125 1552 -91
rect 1506 -163 1552 -125
rect 1506 -197 1512 -163
rect 1546 -197 1552 -163
rect 1506 -235 1552 -197
rect 1506 -269 1512 -235
rect 1546 -269 1552 -235
rect 1506 -307 1552 -269
rect 1506 -341 1512 -307
rect 1546 -341 1552 -307
rect 1506 -379 1552 -341
rect 1506 -413 1512 -379
rect 1546 -413 1552 -379
rect 1506 -451 1552 -413
rect 1506 -485 1512 -451
rect 1546 -485 1552 -451
rect 1506 -523 1552 -485
rect 1506 -557 1512 -523
rect 1546 -557 1552 -523
rect 1506 -600 1552 -557
rect -1496 -647 1496 -641
rect -1496 -681 -1457 -647
rect -1423 -681 -1385 -647
rect -1351 -681 -1313 -647
rect -1279 -681 -1241 -647
rect -1207 -681 -1169 -647
rect -1135 -681 -1097 -647
rect -1063 -681 -1025 -647
rect -991 -681 -953 -647
rect -919 -681 -881 -647
rect -847 -681 -809 -647
rect -775 -681 -737 -647
rect -703 -681 -665 -647
rect -631 -681 -593 -647
rect -559 -681 -521 -647
rect -487 -681 -449 -647
rect -415 -681 -377 -647
rect -343 -681 -305 -647
rect -271 -681 -233 -647
rect -199 -681 -161 -647
rect -127 -681 -89 -647
rect -55 -681 -17 -647
rect 17 -681 55 -647
rect 89 -681 127 -647
rect 161 -681 199 -647
rect 233 -681 271 -647
rect 305 -681 343 -647
rect 377 -681 415 -647
rect 449 -681 487 -647
rect 521 -681 559 -647
rect 593 -681 631 -647
rect 665 -681 703 -647
rect 737 -681 775 -647
rect 809 -681 847 -647
rect 881 -681 919 -647
rect 953 -681 991 -647
rect 1025 -681 1063 -647
rect 1097 -681 1135 -647
rect 1169 -681 1207 -647
rect 1241 -681 1279 -647
rect 1313 -681 1351 -647
rect 1385 -681 1423 -647
rect 1457 -681 1496 -647
rect -1496 -687 1496 -681
<< properties >>
string FIXED_BBOX -1643 -766 1643 766
<< end >>
