magic
tech sky130A
magscale 1 2
timestamp 1731268660
<< nwell >>
rect 24654 16815 26560 16831
rect 24267 15777 26560 16815
rect 25434 14984 26000 15777
<< metal1 >>
rect 22638 17314 22648 17714
rect 23048 17314 23058 17714
<< via1 >>
rect 22648 17314 23048 17714
<< metal2 >>
rect 26209 17839 26308 17849
rect 25135 17789 25234 17799
rect 22648 17714 23048 17724
rect 26209 17732 26308 17742
rect 25135 17682 25234 17692
rect 22648 17304 23048 17314
rect 200 16226 600 16236
rect 600 15826 22386 16226
rect 200 15816 600 15826
rect 22090 2300 22185 15826
rect 27660 4146 27782 4156
rect 27660 4016 27782 4026
rect 25510 3795 25612 3805
rect 25510 3694 25612 3704
rect 25672 2300 25767 3821
rect 25826 3795 25928 3805
rect 25826 3694 25928 3704
rect 22090 2205 25767 2300
<< via2 >>
rect 22648 17314 23048 17714
rect 25135 17692 25234 17789
rect 26209 17742 26308 17839
rect 200 15826 600 16226
rect 27660 4026 27782 4146
rect 25510 3704 25612 3795
rect 25826 3704 25928 3795
<< metal3 >>
rect 26199 17839 26318 17844
rect 25125 17789 25244 17794
rect 22638 17714 23058 17719
rect 22638 17314 22648 17714
rect 23048 17314 23058 17714
rect 25125 17692 25135 17789
rect 25234 17692 25244 17789
rect 26199 17742 26209 17839
rect 26308 17742 26318 17839
rect 26199 17737 26318 17742
rect 25125 17687 25244 17692
rect 22638 17309 23058 17314
rect 190 16226 610 16231
rect 190 15826 200 16226
rect 600 15826 610 16226
rect 190 15821 610 15826
rect 27650 4146 27792 4151
rect 27650 4026 27660 4146
rect 27782 4026 27792 4146
rect 27650 4021 27792 4026
rect 25500 3795 25622 3800
rect 25500 3704 25510 3795
rect 25612 3704 25622 3795
rect 25500 3699 25622 3704
rect 25816 3795 25938 3800
rect 25816 3704 25826 3795
rect 25928 3704 25938 3795
rect 25816 3699 25938 3704
<< via3 >>
rect 22648 17314 23048 17714
rect 25135 17692 25234 17789
rect 26209 17742 26308 17839
rect 200 15826 600 16226
rect 27660 4026 27782 4146
rect 25510 3704 25612 3795
rect 25826 3704 25928 3795
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 200 16227 600 44152
rect 800 17714 1200 44152
rect 18278 18373 18338 45152
rect 18830 18813 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 18830 18753 26289 18813
rect 18278 18313 25214 18373
rect 25154 17790 25214 18313
rect 26229 17840 26289 18753
rect 26208 17839 26309 17840
rect 25134 17789 25235 17790
rect 22647 17714 23049 17715
rect 800 17314 22648 17714
rect 23048 17314 23049 17714
rect 25134 17692 25135 17789
rect 25234 17692 25235 17789
rect 26208 17742 26209 17839
rect 26308 17742 26309 17839
rect 26208 17741 26309 17742
rect 25134 17691 25235 17692
rect 199 16226 601 16227
rect 199 15826 200 16226
rect 600 15826 601 16226
rect 199 15825 601 15826
rect 200 1000 600 15825
rect 800 1000 1200 17314
rect 22647 17313 23049 17314
rect 27659 4146 27783 4147
rect 27659 4026 27660 4146
rect 27782 4105 27783 4146
rect 28766 4105 28826 45152
rect 29318 44952 29378 45152
rect 27782 4045 28826 4105
rect 27782 4026 27783 4045
rect 27659 4025 27783 4026
rect 25470 3795 25650 3854
rect 25470 3704 25510 3795
rect 25612 3704 25650 3795
rect 25470 2706 25650 3704
rect 25789 3795 25969 3851
rect 25789 3704 25826 3795
rect 25928 3704 25969 3795
rect 25789 3082 25969 3704
rect 25789 2902 30542 3082
rect 25470 2526 26678 2706
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 2526
rect 30362 0 30542 2902
use tdc  tdc_0 ~/Documents/Time_Domain_Comparator_ITS/mag
timestamp 1731266514
transform 0 -1 24988 1 0 8540
box -4836 -3709 9311 2246
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 15602 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 15602 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
