* PEX produced on Sen 11 Nov 2024 04:21:00  CST using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from tt_um_tdc_its.ext - technology: sky130A

.subckt tt_um_tdc_its clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6] ua[7]
+ ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0]
+ uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0]
+ uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0]
+ uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] VDPWR VGND
X0 VDPWR.t8 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t3 uo_out[0].t0 VDPWR.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 uo_out[1].t0 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t3 VDPWR.t1 VDPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VGND.t36 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t2 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t6 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t14 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t3 VDPWR.t12 VDPWR.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND.t38 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t2 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t7 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VDPWR.t25 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t4 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t13 VDPWR.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_26743_17057.t0 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t4 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t0 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X7 VDPWR.t36 ua[0].t0 a_25988_7882.t1 VDPWR.t21 sky130_fd_pr__pfet_01v8_lvt ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=15
X8 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t6 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t3 VGND.t10 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_23058_11167.t1 ua[0].t1 VGND.t12 VGND.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=15
X10 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t0 a_25891_11454.t2 a_27981_11167.t0 VGND.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=15
X11 VGND.t43 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t16 a_26743_17057.t1 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X12 VGND.t8 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t4 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t5 VGND.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t15 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t5 VDPWR.t14 VDPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t4 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t6 VGND.t42 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t2 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t5 VGND.t34 VGND.t33 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VDPWR.t27 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t7 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t14 VDPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t2 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t5 VDPWR.t20 VDPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X18 VDPWR.t11 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t6 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t12 VDPWR.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X19 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t1 a_25891_11454.t3 VDPWR.t34 VDPWR.t21 sky130_fd_pr__pfet_01v8_lvt ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=15
X20 a_25914_16928.t0 uo_out[1].t3 VGND.t4 VGND.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X21 VGND.t32 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t7 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t5 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t11 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t8 VDPWR.t35 VDPWR.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t3 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t8 VGND.t19 VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 VGND.t40 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t9 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t2 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 VDPWR.t37 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t9 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t10 VDPWR.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 a_25988_7882.t0 clk.t0 a_25891_11454.t1 VDPWR.t21 sky130_fd_pr__pfet_01v8_lvt ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=15
X27 a_24477_17057.t0 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t4 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t0 VGND.t17 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X28 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t1 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t5 VDPWR.t6 VDPWR.t5 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X29 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t1 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t17 a_26334_16003.t1 VDPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X30 VGND.t15 clk.t1 a_22970_11453.t0 VGND.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=15
X31 a_27981_11167.t1 ua[1].t0 VGND.t44 VGND.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=15
X32 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t9 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t10 VDPWR.t29 VDPWR.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X33 uo_out[1].t1 uo_out[0].t3 a_25456_16928.t1 VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 VDPWR.t33 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t10 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t13 VDPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X35 a_25456_16928.t0 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t6 VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X36 uo_out[0].t1 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t6 a_25914_16928.t1 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X37 VDPWR.t3 ua[1].t1 a_24251_7882.t1 VDPWR.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=15
X38 VGND.t45 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t16 a_24477_17057.t1 VGND.t17 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X39 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t2 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t17 a_24486_16003.t0 VDPWR.t5 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X40 a_26334_16003.t0 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t18 VDPWR.t26 VDPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X41 VGND.t30 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t11 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t15 VGND.t29 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X42 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t12 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t11 VDPWR.t32 VDPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X43 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t1 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t12 VGND.t28 VGND.t27 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X44 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t8 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t13 VDPWR.t10 VDPWR.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X45 VDPWR.t30 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t14 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t7 VDPWR.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X46 VDPWR.t16 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t12 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t11 VDPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X47 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t0 a_22970_11453.t2 a_23058_11167.t0 VGND.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=15
X48 VGND.t26 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t15 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t0 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X49 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t10 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t13 VDPWR.t31 VDPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X50 uo_out[0].t2 uo_out[1].t4 VDPWR.t19 VDPWR.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X51 a_24486_16003.t1 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t18 VDPWR.t17 VDPWR.t5 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X52 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t3 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t16 VGND.t24 VGND.t23 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X53 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t1 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t14 VGND.t6 VGND.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X54 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t1 a_22970_11453.t3 VDPWR.t28 VDPWR.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=15
X55 VGND.t47 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t15 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t0 VGND.t46 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X56 VGND.t14 clk.t2 a_25891_11454.t0 VGND.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=15
X57 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t9 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t16 VDPWR.t22 VDPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X58 VDPWR.t24 uo_out[0].t4 uo_out[1].t2 VDPWR.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X59 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t4 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t17 VGND.t22 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X60 VDPWR.t15 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t17 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t8 VDPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X61 a_24251_7882.t0 clk.t3 a_22970_11453.t1 VDPWR.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=15
R0 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n3 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t5 717.817
R1 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n3 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t4 381.747
R2 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n1 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t3 230.155
R3 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n1 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t6 157.856
R4 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n4 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n1 152
R5 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n0 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t1 99.744
R6 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n2 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t2 84.6561
R7 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n2 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t0 84.0933
R8 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n4 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n0 13.8005
R9 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n0 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n3 8.307
R10 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n0 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n2 6.23388
R11 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n4 4.39453
R12 uo_out[0].n6 uo_out[0].t1 271.209
R13 uo_out[0].n5 uo_out[0].t1 258.846
R14 uo_out[0].n1 uo_out[0].t4 230.155
R15 uo_out[0].n3 uo_out[0].n0 193.548
R16 uo_out[0].n1 uo_out[0].t3 157.856
R17 uo_out[0].n2 uo_out[0].n1 152
R18 uo_out[0].n7 uo_out[0] 33.8304
R19 uo_out[0] uo_out[0].n3 31.2308
R20 uo_out[0].n0 uo_out[0].t0 26.5955
R21 uo_out[0].n0 uo_out[0].t2 26.5955
R22 uo_out[0].n3 uo_out[0].n2 23.8989
R23 uo_out[0] uo_out[0].n6 14.2478
R24 uo_out[0].n2 uo_out[0] 4.39453
R25 uo_out[0].n4 uo_out[0] 3.76521
R26 uo_out[0].n5 uo_out[0].n4 3.03935
R27 uo_out[0] uo_out[0].n5 2.30266
R28 uo_out[0].n7 uo_out[0] 1.80364
R29 uo_out[0].n4 uo_out[0] 0.921363
R30 uo_out[0].n6 uo_out[0] 0.829277
R31 uo_out[0] uo_out[0].n7 0.00555051
R32 VDPWR.n170 VDPWR.n8 8442.35
R33 VDPWR.n170 VDPWR.n6 8442.35
R34 VDPWR.n169 VDPWR.n15 8442.35
R35 VDPWR.n169 VDPWR.n16 8442.35
R36 VDPWR.n152 VDPWR.n142 8442.35
R37 VDPWR.n152 VDPWR.n139 8442.35
R38 VDPWR.n26 VDPWR.n25 8442.35
R39 VDPWR.n26 VDPWR.n18 8442.35
R40 VDPWR.n161 VDPWR.n8 5738.82
R41 VDPWR.n14 VDPWR.n4 5738.82
R42 VDPWR.n11 VDPWR.n4 5738.82
R43 VDPWR.n11 VDPWR.n6 5738.82
R44 VDPWR.n15 VDPWR.n14 5738.82
R45 VDPWR.n160 VDPWR.n16 5738.82
R46 VDPWR.n162 VDPWR.n160 5738.82
R47 VDPWR.n162 VDPWR.n161 5738.82
R48 VDPWR.n142 VDPWR.n141 5738.82
R49 VDPWR.n145 VDPWR.n21 5738.82
R50 VDPWR.n145 VDPWR.n144 5738.82
R51 VDPWR.n144 VDPWR.n139 5738.82
R52 VDPWR.n25 VDPWR.n21 5738.82
R53 VDPWR.n22 VDPWR.n18 5738.82
R54 VDPWR.n140 VDPWR.n22 5738.82
R55 VDPWR.n141 VDPWR.n140 5738.82
R56 VDPWR.n12 VDPWR.n11 2703.53
R57 VDPWR.n161 VDPWR.n12 2703.53
R58 VDPWR.n14 VDPWR.n13 2703.53
R59 VDPWR.n160 VDPWR.n13 2703.53
R60 VDPWR.n144 VDPWR.n27 2703.53
R61 VDPWR.n141 VDPWR.n27 2703.53
R62 VDPWR.n153 VDPWR.n21 2703.53
R63 VDPWR.n153 VDPWR.n22 2703.53
R64 VDPWR.n119 VDPWR.n37 2142.35
R65 VDPWR.n37 VDPWR.n29 2142.35
R66 VDPWR.n135 VDPWR.n30 2142.35
R67 VDPWR.n125 VDPWR.n30 2142.35
R68 VDPWR.n111 VDPWR.n86 2142.35
R69 VDPWR.n111 VDPWR.n85 2142.35
R70 VDPWR.n110 VDPWR.n91 2142.35
R71 VDPWR.n110 VDPWR.n92 2142.35
R72 VDPWR.n129 VDPWR.n36 1644.71
R73 VDPWR.n129 VDPWR.n128 1644.71
R74 VDPWR.n120 VDPWR.n31 1644.71
R75 VDPWR.n121 VDPWR.n120 1644.71
R76 VDPWR.n102 VDPWR.n89 1644.71
R77 VDPWR.n95 VDPWR.n89 1644.71
R78 VDPWR.n101 VDPWR.n90 1644.71
R79 VDPWR.n94 VDPWR.n90 1644.71
R80 VDPWR.n171 VDPWR.n7 752.211
R81 VDPWR.n168 VDPWR.n167 752.211
R82 VDPWR.n151 VDPWR.n143 752.211
R83 VDPWR.n24 VDPWR.n17 752.211
R84 VDPWR.n159 VDPWR.n7 612.141
R85 VDPWR.n167 VDPWR.n166 612.141
R86 VDPWR.n166 VDPWR.n163 612.141
R87 VDPWR.n163 VDPWR.n159 612.141
R88 VDPWR.n147 VDPWR.n143 612.141
R89 VDPWR.n146 VDPWR.n19 612.141
R90 VDPWR.n147 VDPWR.n146 612.141
R91 VDPWR.n24 VDPWR.n19 612.141
R92 VDPWR.n128 VDPWR.n119 497.647
R93 VDPWR.n31 VDPWR.n28 497.647
R94 VDPWR.n36 VDPWR.n28 497.647
R95 VDPWR.n36 VDPWR.n29 497.647
R96 VDPWR.n135 VDPWR.n31 497.647
R97 VDPWR.n125 VDPWR.n121 497.647
R98 VDPWR.n127 VDPWR.n121 497.647
R99 VDPWR.n128 VDPWR.n127 497.647
R100 VDPWR.n95 VDPWR.n86 497.647
R101 VDPWR.n103 VDPWR.n101 497.647
R102 VDPWR.n103 VDPWR.n102 497.647
R103 VDPWR.n102 VDPWR.n85 497.647
R104 VDPWR.n101 VDPWR.n91 497.647
R105 VDPWR.n94 VDPWR.n92 497.647
R106 VDPWR.n96 VDPWR.n94 497.647
R107 VDPWR.n96 VDPWR.n95 497.647
R108 VDPWR.n172 VDPWR.n171 440.687
R109 VDPWR.n168 VDPWR.n158 440.687
R110 VDPWR.n151 VDPWR.n150 440.687
R111 VDPWR.n156 VDPWR.n17 440.687
R112 VDPWR.t4 VDPWR.n87 420.019
R113 VDPWR.t4 VDPWR.n88 420.019
R114 VDPWR.n136 VDPWR.t5 420.019
R115 VDPWR.n126 VDPWR.t5 420.019
R116 VDPWR.n61 VDPWR.t11 342.377
R117 VDPWR.n61 VDPWR.t33 342.375
R118 VDPWR.n49 VDPWR.t29 338.892
R119 VDPWR.n49 VDPWR.t31 338.892
R120 VDPWR.n42 VDPWR.n40 327.377
R121 VDPWR.n55 VDPWR.n43 327.377
R122 VDPWR.n47 VDPWR.n45 327.377
R123 VDPWR.n42 VDPWR.n41 327.375
R124 VDPWR.n55 VDPWR.n44 327.375
R125 VDPWR.n47 VDPWR.n46 327.375
R126 VDPWR.n158 VDPWR.n3 300.435
R127 VDPWR.n174 VDPWR.n3 300.435
R128 VDPWR.n174 VDPWR.n173 300.435
R129 VDPWR.n173 VDPWR.n172 300.435
R130 VDPWR.n156 VDPWR.n155 300.435
R131 VDPWR.n155 VDPWR.n1 300.435
R132 VDPWR.n149 VDPWR.n1 300.435
R133 VDPWR.n150 VDPWR.n149 300.435
R134 VDPWR.n159 VDPWR.n5 288.377
R135 VDPWR.n166 VDPWR.n165 288.377
R136 VDPWR.n148 VDPWR.n147 288.377
R137 VDPWR.n154 VDPWR.n19 288.377
R138 VDPWR.n173 VDPWR.n5 281.976
R139 VDPWR.n165 VDPWR.n3 281.976
R140 VDPWR.n149 VDPWR.n148 281.976
R141 VDPWR.n155 VDPWR.n154 281.976
R142 VDPWR.n73 VDPWR.t24 249.362
R143 VDPWR.n65 VDPWR.t8 249.362
R144 VDPWR.n75 VDPWR.t1 247.394
R145 VDPWR.n68 VDPWR.t19 247.394
R146 VDPWR.n134 VDPWR.n32 228.518
R147 VDPWR.n124 VDPWR.n32 228.518
R148 VDPWR.n117 VDPWR.n34 228.518
R149 VDPWR.n118 VDPWR.n117 228.518
R150 VDPWR.n112 VDPWR.n84 228.518
R151 VDPWR.n112 VDPWR.n83 228.518
R152 VDPWR.n109 VDPWR.n93 228.518
R153 VDPWR.n109 VDPWR.n108 228.518
R154 VDPWR.n133 VDPWR.n33 175.435
R155 VDPWR.n123 VDPWR.n33 175.435
R156 VDPWR.n131 VDPWR.n130 175.435
R157 VDPWR.n130 VDPWR.n35 175.435
R158 VDPWR.n100 VDPWR.n99 175.435
R159 VDPWR.n99 VDPWR.n98 175.435
R160 VDPWR.n106 VDPWR.n105 175.435
R161 VDPWR.n107 VDPWR.n106 175.435
R162 VDPWR.n137 VDPWR.t23 173.055
R163 VDPWR.n88 VDPWR.t7 166.746
R164 VDPWR.n137 VDPWR.t9 123.913
R165 VDPWR VDPWR.t13 109.584
R166 VDPWR VDPWR.n136 107.258
R167 VDPWR.n137 VDPWR 100.95
R168 VDPWR.n108 VDPWR.n92 92.5005
R169 VDPWR.n92 VDPWR.n88 92.5005
R170 VDPWR.n97 VDPWR.n96 92.5005
R171 VDPWR.n96 VDPWR.n88 92.5005
R172 VDPWR.n86 VDPWR.n84 92.5005
R173 VDPWR.n88 VDPWR.n86 92.5005
R174 VDPWR.n85 VDPWR.n83 92.5005
R175 VDPWR.n87 VDPWR.n85 92.5005
R176 VDPWR.n104 VDPWR.n103 92.5005
R177 VDPWR.n103 VDPWR.n87 92.5005
R178 VDPWR.n93 VDPWR.n91 92.5005
R179 VDPWR.n91 VDPWR.n87 92.5005
R180 VDPWR.n125 VDPWR.n124 92.5005
R181 VDPWR.n126 VDPWR.n125 92.5005
R182 VDPWR.n127 VDPWR.n122 92.5005
R183 VDPWR.n127 VDPWR.n126 92.5005
R184 VDPWR.n119 VDPWR.n118 92.5005
R185 VDPWR.n126 VDPWR.n119 92.5005
R186 VDPWR.n34 VDPWR.n29 92.5005
R187 VDPWR.n136 VDPWR.n29 92.5005
R188 VDPWR.n132 VDPWR.n28 92.5005
R189 VDPWR.n136 VDPWR.n28 92.5005
R190 VDPWR.n135 VDPWR.n134 92.5005
R191 VDPWR.n136 VDPWR.n135 92.5005
R192 VDPWR.n78 VDPWR.t6 89.8482
R193 VDPWR.n81 VDPWR.t20 89.8122
R194 VDPWR.n116 VDPWR.t17 84.664
R195 VDPWR.n113 VDPWR.t26 84.664
R196 VDPWR.t7 VDPWR.t18 75.7121
R197 VDPWR.t23 VDPWR.t0 75.7121
R198 VDPWR.t21 VDPWR.n23 73.0334
R199 VDPWR.t21 VDPWR.n138 73.0334
R200 VDPWR.t2 VDPWR.n9 73.0334
R201 VDPWR.t2 VDPWR.n10 73.0334
R202 VDPWR.t18 VDPWR 63.0935
R203 VDPWR.t0 VDPWR 63.0935
R204 VDPWR.n134 VDPWR.n133 53.0829
R205 VDPWR.n124 VDPWR.n123 53.0829
R206 VDPWR.n123 VDPWR.n122 53.0829
R207 VDPWR.n122 VDPWR.n35 53.0829
R208 VDPWR.n133 VDPWR.n132 53.0829
R209 VDPWR.n132 VDPWR.n131 53.0829
R210 VDPWR.n131 VDPWR.n34 53.0829
R211 VDPWR.n118 VDPWR.n35 53.0829
R212 VDPWR.n98 VDPWR.n84 53.0829
R213 VDPWR.n105 VDPWR.n104 53.0829
R214 VDPWR.n104 VDPWR.n100 53.0829
R215 VDPWR.n100 VDPWR.n83 53.0829
R216 VDPWR.n105 VDPWR.n93 53.0829
R217 VDPWR.n108 VDPWR.n107 53.0829
R218 VDPWR.n107 VDPWR.n97 53.0829
R219 VDPWR.n98 VDPWR.n97 53.0829
R220 VDPWR.n164 VDPWR.t28 39.7543
R221 VDPWR.n164 VDPWR.t3 39.7543
R222 VDPWR.n20 VDPWR.t34 39.7543
R223 VDPWR.n20 VDPWR.t36 39.7543
R224 VDPWR.n60 VDPWR.n38 34.6358
R225 VDPWR.n50 VDPWR.n47 31.624
R226 VDPWR.n56 VDPWR.n55 30.8711
R227 VDPWR.n41 VDPWR.t22 26.5955
R228 VDPWR.n41 VDPWR.t15 26.5955
R229 VDPWR.n40 VDPWR.t10 26.5955
R230 VDPWR.n40 VDPWR.t30 26.5955
R231 VDPWR.n44 VDPWR.t14 26.5955
R232 VDPWR.n44 VDPWR.t27 26.5955
R233 VDPWR.n43 VDPWR.t12 26.5955
R234 VDPWR.n43 VDPWR.t25 26.5955
R235 VDPWR.n46 VDPWR.t32 26.5955
R236 VDPWR.n46 VDPWR.t16 26.5955
R237 VDPWR.n45 VDPWR.t35 26.5955
R238 VDPWR.n45 VDPWR.t37 26.5955
R239 VDPWR.n74 VDPWR.n73 25.977
R240 VDPWR.n67 VDPWR.n65 25.977
R241 VDPWR.n55 VDPWR.n54 25.6005
R242 VDPWR.n54 VDPWR.n47 24.8476
R243 VDPWR.n75 VDPWR.n74 24.4711
R244 VDPWR.n68 VDPWR.n67 24.4711
R245 VDPWR.n56 VDPWR.n42 19.577
R246 VDPWR.n50 VDPWR.n49 18.824
R247 VDPWR.n106 VDPWR.n90 16.8187
R248 VDPWR.t4 VDPWR.n90 16.8187
R249 VDPWR.n99 VDPWR.n89 16.8187
R250 VDPWR.t4 VDPWR.n89 16.8187
R251 VDPWR.n112 VDPWR.n111 16.8187
R252 VDPWR.n111 VDPWR.t4 16.8187
R253 VDPWR.n110 VDPWR.n109 16.8187
R254 VDPWR.t4 VDPWR.n110 16.8187
R255 VDPWR.n120 VDPWR.n33 16.8187
R256 VDPWR.n120 VDPWR.t5 16.8187
R257 VDPWR.n130 VDPWR.n129 16.8187
R258 VDPWR.n129 VDPWR.t5 16.8187
R259 VDPWR.n117 VDPWR.n37 16.8187
R260 VDPWR.n37 VDPWR.t5 16.8187
R261 VDPWR.n32 VDPWR.n30 16.8187
R262 VDPWR.n30 VDPWR.t5 16.8187
R263 VDPWR.n137 VDPWR 14.3306
R264 VDPWR.n61 VDPWR.n60 13.5534
R265 VDPWR.n62 VDPWR.n61 11.1829
R266 VDPWR.n138 VDPWR.n137 10.0115
R267 VDPWR.n137 VDPWR.n9 9.53482
R268 VDPWR.n49 VDPWR.n48 9.3005
R269 VDPWR.n51 VDPWR.n50 9.3005
R270 VDPWR.n52 VDPWR.n47 9.3005
R271 VDPWR.n54 VDPWR.n53 9.3005
R272 VDPWR.n55 VDPWR.n39 9.3005
R273 VDPWR.n57 VDPWR.n56 9.3005
R274 VDPWR.n58 VDPWR.n38 9.3005
R275 VDPWR.n60 VDPWR.n59 9.3005
R276 VDPWR.n69 VDPWR.n68 9.3005
R277 VDPWR.n65 VDPWR.n63 9.3005
R278 VDPWR.n67 VDPWR.n66 9.3005
R279 VDPWR.n76 VDPWR.n75 9.3005
R280 VDPWR.n73 VDPWR.n72 9.3005
R281 VDPWR.n74 VDPWR.n71 9.3005
R282 VDPWR.n165 VDPWR.n13 9.2505
R283 VDPWR.t2 VDPWR.n13 9.2505
R284 VDPWR.n12 VDPWR.n5 9.2505
R285 VDPWR.t2 VDPWR.n12 9.2505
R286 VDPWR.n171 VDPWR.n170 9.2505
R287 VDPWR.n170 VDPWR.t2 9.2505
R288 VDPWR.n169 VDPWR.n168 9.2505
R289 VDPWR.t2 VDPWR.n169 9.2505
R290 VDPWR.n152 VDPWR.n151 9.2505
R291 VDPWR.t21 VDPWR.n152 9.2505
R292 VDPWR.n148 VDPWR.n27 9.2505
R293 VDPWR.t21 VDPWR.n27 9.2505
R294 VDPWR.n154 VDPWR.n153 9.2505
R295 VDPWR.n153 VDPWR.t21 9.2505
R296 VDPWR.n26 VDPWR.n17 9.2505
R297 VDPWR.t21 VDPWR.n26 9.2505
R298 VDPWR VDPWR.n176 6.23715
R299 VDPWR.n79 VDPWR.n70 4.51973
R300 VDPWR.n80 VDPWR.n64 4.51973
R301 VDPWR.n82 VDPWR.n81 4.51973
R302 VDPWR.n78 VDPWR.n77 4.51973
R303 VDPWR.n167 VDPWR.n16 4.02224
R304 VDPWR.n16 VDPWR.n10 4.02224
R305 VDPWR.n163 VDPWR.n162 4.02224
R306 VDPWR.n162 VDPWR.n10 4.02224
R307 VDPWR.n8 VDPWR.n7 4.02224
R308 VDPWR.n10 VDPWR.n8 4.02224
R309 VDPWR.n172 VDPWR.n6 4.02224
R310 VDPWR.n9 VDPWR.n6 4.02224
R311 VDPWR.n174 VDPWR.n4 4.02224
R312 VDPWR.n9 VDPWR.n4 4.02224
R313 VDPWR.n158 VDPWR.n15 4.02224
R314 VDPWR.n15 VDPWR.n9 4.02224
R315 VDPWR.n146 VDPWR.n145 4.02224
R316 VDPWR.n145 VDPWR.n23 4.02224
R317 VDPWR.n143 VDPWR.n139 4.02224
R318 VDPWR.n139 VDPWR.n23 4.02224
R319 VDPWR.n25 VDPWR.n24 4.02224
R320 VDPWR.n25 VDPWR.n23 4.02224
R321 VDPWR.n156 VDPWR.n18 4.02224
R322 VDPWR.n138 VDPWR.n18 4.02224
R323 VDPWR.n140 VDPWR.n1 4.02224
R324 VDPWR.n140 VDPWR.n138 4.02224
R325 VDPWR.n150 VDPWR.n142 4.02224
R326 VDPWR.n142 VDPWR.n138 4.02224
R327 VDPWR.n175 VDPWR.n2 2.29309
R328 VDPWR.n42 VDPWR.n38 2.25932
R329 VDPWR.n157 VDPWR 1.28325
R330 VDPWR.n114 VDPWR.n82 1.27487
R331 VDPWR.n2 VDPWR 1.2145
R332 VDPWR.n117 VDPWR.n116 1.20034
R333 VDPWR.n113 VDPWR.n112 1.20034
R334 VDPWR.n157 VDPWR.n0 1.12277
R335 VDPWR.n116 VDPWR.n115 0.771119
R336 VDPWR.n176 VDPWR.n0 0.708833
R337 VDPWR.n80 VDPWR.n79 0.663962
R338 VDPWR.n165 VDPWR.n164 0.489974
R339 VDPWR.n154 VDPWR.n20 0.489974
R340 VDPWR.n79 VDPWR.n78 0.445212
R341 VDPWR.n81 VDPWR.n80 0.442808
R342 VDPWR.n176 VDPWR.n175 0.414434
R343 VDPWR.n114 VDPWR.n113 0.405139
R344 VDPWR.n164 VDPWR.n0 0.40437
R345 VDPWR.n20 VDPWR.n0 0.40437
R346 VDPWR.n115 VDPWR.n114 0.343284
R347 VDPWR.n70 VDPWR 0.28826
R348 VDPWR VDPWR.n62 0.278625
R349 VDPWR.n150 VDPWR.n2 0.216779
R350 VDPWR.n172 VDPWR.n2 0.216779
R351 VDPWR.n157 VDPWR.n156 0.216779
R352 VDPWR.n175 VDPWR.n1 0.216779
R353 VDPWR.n158 VDPWR.n157 0.216779
R354 VDPWR.n175 VDPWR.n174 0.216779
R355 VDPWR.n66 VDPWR.n63 0.120292
R356 VDPWR.n72 VDPWR.n71 0.120292
R357 VDPWR.n77 VDPWR.n71 0.112479
R358 VDPWR.n66 VDPWR.n64 0.108573
R359 VDPWR.n59 VDPWR.n58 0.0963333
R360 VDPWR.n58 VDPWR.n57 0.0963333
R361 VDPWR.n57 VDPWR.n39 0.0963333
R362 VDPWR.n53 VDPWR.n39 0.0963333
R363 VDPWR.n53 VDPWR.n52 0.0963333
R364 VDPWR.n52 VDPWR.n51 0.0963333
R365 VDPWR.n51 VDPWR.n48 0.0963333
R366 VDPWR.n59 VDPWR 0.078625
R367 VDPWR.n115 VDPWR 0.0505
R368 VDPWR.n48 VDPWR 0.0484167
R369 VDPWR VDPWR.n69 0.0239375
R370 VDPWR.n76 VDPWR 0.0239375
R371 VDPWR.n62 VDPWR 0.0182083
R372 VDPWR.n82 VDPWR.n63 0.0122188
R373 VDPWR.n69 VDPWR.n64 0.0122188
R374 VDPWR.n72 VDPWR.n70 0.00961458
R375 VDPWR.n77 VDPWR.n76 0.0083125
R376 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n2 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t5 717.539
R377 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n2 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t4 382.024
R378 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n1 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t3 229.369
R379 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n1 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t6 157.07
R380 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n4 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n1 152
R381 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n0 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t2 99.4459
R382 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n3 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t0 84.4033
R383 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n3 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t1 84.3461
R384 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n4 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n0 13.9367
R385 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n0 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n2 8.31548
R386 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n0 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n3 6.2204
R387 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n4 5.92643
R388 uo_out[1].n5 uo_out[1].t1 271.209
R389 uo_out[1].n4 uo_out[1].t1 258.846
R390 uo_out[1].n0 uo_out[1].t4 229.369
R391 uo_out[1] uo_out[1].n2 224.778
R392 uo_out[1].n0 uo_out[1].t3 157.07
R393 uo_out[1].n1 uo_out[1].n0 152
R394 uo_out[1].n7 uo_out[1] 33.4599
R395 uo_out[1].n2 uo_out[1].t2 26.5955
R396 uo_out[1].n2 uo_out[1].t0 26.5955
R397 uo_out[1].n6 uo_out[1].n1 10.0773
R398 uo_out[1].n6 uo_out[1].n5 9.3005
R399 uo_out[1].n1 uo_out[1] 5.92643
R400 uo_out[1] uo_out[1].n6 5.41118
R401 uo_out[1].n3 uo_out[1] 3.76521
R402 uo_out[1].n4 uo_out[1].n3 3.03935
R403 uo_out[1] uo_out[1].n4 2.30266
R404 uo_out[1].n7 uo_out[1] 1.68191
R405 uo_out[1].n3 uo_out[1] 0.921363
R406 uo_out[1].n5 uo_out[1] 0.829277
R407 uo_out[1] uo_out[1].n7 0.0712071
R408 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n14 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t10 212.081
R409 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n13 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t9 212.081
R410 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n1 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t8 212.081
R411 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n10 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t4 212.081
R412 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n2 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t3 212.081
R413 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n7 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t14 212.081
R414 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n5 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t13 212.081
R415 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n3 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t6 212.081
R416 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n4 tdc_0.sky130_fd_sc_hd__inv_8_0.A 171.969
R417 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n6 tdc_0.sky130_fd_sc_hd__inv_8_0.A 152
R418 tdc_0.sky130_fd_sc_hd__inv_8_0.A tdc_0.sky130_fd_sc_hd__inv_8_0.A.n8 152
R419 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n9 tdc_0.sky130_fd_sc_hd__inv_8_0.A 152
R420 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n0 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n11 152
R421 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n12 tdc_0.sky130_fd_sc_hd__inv_8_0.A 152
R422 tdc_0.sky130_fd_sc_hd__inv_8_0.A tdc_0.sky130_fd_sc_hd__inv_8_0.A.n15 152
R423 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n14 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t16 139.78
R424 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n13 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t15 139.78
R425 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n1 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t12 139.78
R426 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n10 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t7 139.78
R427 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n2 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t5 139.78
R428 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n7 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t2 139.78
R429 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n5 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t17 139.78
R430 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n3 tdc_0.sky130_fd_sc_hd__inv_8_0.A.t11 139.78
R431 tdc_0.sky130_fd_sc_hd__inv_8_0.A tdc_0.sky130_fd_sc_hd__inv_8_0.A.n0 43.0085
R432 tdc_0.sky130_fd_sc_hd__inv_8_0.A tdc_0.sky130_fd_sc_hd__inv_8_0.A.t0 42.6438
R433 tdc_0.sky130_fd_sc_hd__inv_8_0.A tdc_0.sky130_fd_sc_hd__inv_8_0.A.t1 39.7543
R434 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n4 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n3 30.6732
R435 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n5 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n4 30.6732
R436 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n6 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n5 30.6732
R437 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n7 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n6 30.6732
R438 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n8 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n7 30.6732
R439 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n8 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n2 30.6732
R440 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n9 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n2 30.6732
R441 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n10 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n9 30.6732
R442 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n11 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n10 30.6732
R443 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n11 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n1 30.6732
R444 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n12 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n1 30.6732
R445 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n13 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n12 30.6732
R446 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n15 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n13 30.6732
R447 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n15 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n14 30.6732
R448 tdc_0.sky130_fd_sc_hd__inv_8_0.A.n0 tdc_0.sky130_fd_sc_hd__inv_8_0.A 26.6304
R449 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t17 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t16 1119.58
R450 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n0 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t17 731.562
R451 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n0 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t18 723.615
R452 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t18 tdc_0.sky130_fd_sc_hd__inv_8_0.Y 721.894
R453 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n14 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n3 205.28
R454 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n13 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n4 205.28
R455 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n17 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n2 205.28
R456 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n16 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n15 205.28
R457 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n12 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n5 99.1759
R458 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n11 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n6 99.1759
R459 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n10 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n7 99.1759
R460 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n9 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n8 99.1759
R461 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n14 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n13 38.4005
R462 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n17 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n16 38.4005
R463 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n16 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n14 38.4005
R464 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n12 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n11 34.3584
R465 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n11 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n10 34.3584
R466 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n10 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n9 34.3584
R467 tdc_0.sky130_fd_sc_hd__inv_8_0.Y tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n12 32.411
R468 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n9 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n1 30.9412
R469 tdc_0.sky130_fd_sc_hd__inv_8_0.Y tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n17 30.14
R470 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n13 tdc_0.sky130_fd_sc_hd__inv_8_0.Y 27.6358
R471 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n3 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t13 26.5955
R472 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n3 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t11 26.5955
R473 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n4 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t10 26.5955
R474 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n4 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t9 26.5955
R475 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n2 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t12 26.5955
R476 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n2 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t8 26.5955
R477 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n15 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t7 26.5955
R478 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n15 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t14 26.5955
R479 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n5 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t0 24.9236
R480 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n5 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t3 24.9236
R481 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n6 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t5 24.9236
R482 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n6 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t1 24.9236
R483 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n7 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t6 24.9236
R484 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n7 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t2 24.9236
R485 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n8 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t15 24.9236
R486 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n8 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t4 24.9236
R487 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n1 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n0 15.1977
R488 tdc_0.sky130_fd_sc_hd__inv_8_0.Y tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n1 3.15412
R489 VGND.n137 VGND.n136 177953
R490 VGND.n119 VGND.n27 177460
R491 VGND.n27 VGND.n26 24287.8
R492 VGND.n149 VGND.n141 11489.7
R493 VGND.n141 VGND.n28 11489.7
R494 VGND.n87 VGND.n80 11489.7
R495 VGND.n80 VGND.n76 11489.7
R496 VGND.n97 VGND.n82 11489.7
R497 VGND.n97 VGND.n83 11489.7
R498 VGND.n155 VGND.n29 11489.7
R499 VGND.n151 VGND.n29 11489.7
R500 VGND.n149 VGND.n140 9421.24
R501 VGND.n87 VGND.n77 9421.24
R502 VGND.n100 VGND.n75 9421.24
R503 VGND.n100 VGND.n99 9421.24
R504 VGND.n99 VGND.n76 9421.24
R505 VGND.n82 VGND.n75 9421.24
R506 VGND.n90 VGND.n83 9421.24
R507 VGND.n91 VGND.n90 9421.24
R508 VGND.n91 VGND.n77 9421.24
R509 VGND.n155 VGND.n24 9421.24
R510 VGND.n151 VGND.n33 9421.24
R511 VGND.n139 VGND.n33 9421.24
R512 VGND.n140 VGND.n139 9421.24
R513 VGND.n157 VGND.n24 9421.24
R514 VGND.n157 VGND.n25 9421.24
R515 VGND.n28 VGND.n25 9421.24
R516 VGND.n150 VGND.n138 4765.62
R517 VGND.n156 VGND.n27 3476.72
R518 VGND.n116 VGND.n46 2306.06
R519 VGND.n120 VGND.n116 2306.06
R520 VGND.n126 VGND.n47 2306.06
R521 VGND.n115 VGND.n47 2306.06
R522 VGND.n43 VGND.n35 2306.06
R523 VGND.n129 VGND.n43 2306.06
R524 VGND.n135 VGND.n36 2306.06
R525 VGND.n42 VGND.n36 2306.06
R526 VGND.n99 VGND.n98 2068.5
R527 VGND.n98 VGND.n77 2068.5
R528 VGND.n81 VGND.n75 2068.5
R529 VGND.n90 VGND.n81 2068.5
R530 VGND.n33 VGND.n32 2068.5
R531 VGND.n32 VGND.n24 2068.5
R532 VGND.n143 VGND.n140 2068.5
R533 VGND.n143 VGND.n25 2068.5
R534 VGND.n122 VGND.n48 1489.09
R535 VGND.n122 VGND.n121 1489.09
R536 VGND.n131 VGND.n37 1489.09
R537 VGND.n131 VGND.n130 1489.09
R538 VGND.n48 VGND.n46 816.971
R539 VGND.n126 VGND.n48 816.971
R540 VGND.n121 VGND.n115 816.971
R541 VGND.n121 VGND.n120 816.971
R542 VGND.n37 VGND.n35 816.971
R543 VGND.n135 VGND.n37 816.971
R544 VGND.n130 VGND.n42 816.971
R545 VGND.n130 VGND.n129 816.971
R546 VGND.n138 VGND.n137 730.953
R547 VGND.n88 VGND.n86 677.422
R548 VGND.n96 VGND.n95 677.422
R549 VGND.n153 VGND.n152 677.422
R550 VGND.n148 VGND.n147 677.422
R551 VGND.n89 VGND.n88 612.141
R552 VGND.n95 VGND.n94 612.141
R553 VGND.n94 VGND.n92 612.141
R554 VGND.n92 VGND.n89 612.141
R555 VGND.n142 VGND.n30 612.141
R556 VGND.n145 VGND.n142 612.141
R557 VGND.n152 VGND.n30 612.141
R558 VGND.n148 VGND.n145 612.141
R559 VGND.t21 VGND.t29 320.555
R560 VGND.t35 VGND.t21 320.555
R561 VGND.t33 VGND.t31 320.555
R562 VGND.t31 VGND.t27 320.555
R563 VGND.t27 VGND.t25 320.555
R564 VGND.t25 VGND.t23 320.555
R565 VGND.t18 VGND.t37 316.711
R566 VGND.t39 VGND.t18 316.711
R567 VGND.t5 VGND.t46 316.711
R568 VGND.t46 VGND.t9 316.711
R569 VGND.t9 VGND.t7 316.711
R570 VGND.t7 VGND.t41 316.711
R571 VGND.n42 VGND.n41 292.5
R572 VGND.n128 VGND.n42 292.5
R573 VGND.n129 VGND.n45 292.5
R574 VGND.n129 VGND.n128 292.5
R575 VGND.n39 VGND.n35 292.5
R576 VGND.n136 VGND.n35 292.5
R577 VGND.n135 VGND.n134 292.5
R578 VGND.n136 VGND.n135 292.5
R579 VGND.n115 VGND.n114 292.5
R580 VGND.n119 VGND.n115 292.5
R581 VGND.n120 VGND.n118 292.5
R582 VGND.n120 VGND.n119 292.5
R583 VGND.n112 VGND.n46 292.5
R584 VGND.n127 VGND.n46 292.5
R585 VGND.n126 VGND.n125 292.5
R586 VGND.n127 VGND.n126 292.5
R587 VGND.n69 VGND.t30 291.606
R588 VGND.n19 VGND.t38 291.606
R589 VGND.n56 VGND.t24 284.024
R590 VGND.n6 VGND.t42 284.024
R591 VGND.t29 VGND 244.232
R592 VGND.t37 VGND 241.303
R593 VGND.n60 VGND.n55 213.613
R594 VGND.n53 VGND.n52 213.613
R595 VGND.n67 VGND.n66 213.613
R596 VGND.n10 VGND.n5 213.613
R597 VGND.n3 VGND.n2 213.613
R598 VGND.n17 VGND.n16 213.613
R599 VGND.n138 VGND.n34 192.534
R600 VGND.n86 VGND.n85 187.236
R601 VGND.n96 VGND.n84 187.236
R602 VGND.n154 VGND.n153 187.236
R603 VGND.n147 VGND.n146 187.236
R604 VGND.n137 VGND.t35 183.174
R605 VGND.n26 VGND.t39 180.977
R606 VGND.n50 VGND.t4 157.988
R607 VGND.n49 VGND.t1 157.988
R608 VGND.t13 VGND.n34 157.649
R609 VGND.t13 VGND.n79 157.649
R610 VGND.n117 VGND.n112 149.835
R611 VGND.n118 VGND.n117 149.835
R612 VGND.n114 VGND.n111 149.835
R613 VGND.n125 VGND.n111 149.835
R614 VGND.n44 VGND.n39 149.835
R615 VGND.n45 VGND.n44 149.835
R616 VGND.n41 VGND.n38 149.835
R617 VGND.n134 VGND.n38 149.835
R618 VGND.n137 VGND.t33 137.381
R619 VGND.n26 VGND.t5 135.733
R620 VGND.n89 VGND.n78 134.4
R621 VGND.n94 VGND.n93 134.4
R622 VGND.n31 VGND.n30 134.4
R623 VGND.n145 VGND.n144 134.4
R624 VGND.n78 VGND.n74 128
R625 VGND.n93 VGND.n73 128
R626 VGND.n31 VGND.n22 128
R627 VGND.n144 VGND.n23 128
R628 VGND.n84 VGND.n73 123.709
R629 VGND.n101 VGND.n74 123.709
R630 VGND.n85 VGND.n74 123.709
R631 VGND.n154 VGND.n22 123.709
R632 VGND.n158 VGND.n23 123.709
R633 VGND.n146 VGND.n23 123.709
R634 VGND.n102 VGND.n73 122.353
R635 VGND.n159 VGND.n22 122.353
R636 VGND.n132 VGND.n131 117.001
R637 VGND.n131 VGND.t2 117.001
R638 VGND.n44 VGND.n43 117.001
R639 VGND.n43 VGND.t2 117.001
R640 VGND.n38 VGND.n36 117.001
R641 VGND.n36 VGND.t2 117.001
R642 VGND.n123 VGND.n122 117.001
R643 VGND.n122 VGND.t17 117.001
R644 VGND.n117 VGND.n116 117.001
R645 VGND.n116 VGND.t17 117.001
R646 VGND.n111 VGND.n47 117.001
R647 VGND.n47 VGND.t17 117.001
R648 VGND.n150 VGND.t11 107.222
R649 VGND.n156 VGND.t11 107.222
R650 VGND.n124 VGND.n123 96.7534
R651 VGND.n123 VGND.n113 96.7534
R652 VGND.n133 VGND.n132 96.7534
R653 VGND.n132 VGND.n40 96.7534
R654 VGND.n128 VGND.t16 93.7267
R655 VGND.n108 VGND.t45 84.028
R656 VGND.n106 VGND.t43 84.028
R657 VGND VGND.n127 83.4681
R658 VGND.n93 VGND.n81 73.1255
R659 VGND.t13 VGND.n81 73.1255
R660 VGND.n98 VGND.n78 73.1255
R661 VGND.n98 VGND.t13 73.1255
R662 VGND.n86 VGND.n80 73.1255
R663 VGND.t13 VGND.n80 73.1255
R664 VGND.n97 VGND.n96 73.1255
R665 VGND.t13 VGND.n97 73.1255
R666 VGND.n153 VGND.n29 73.1255
R667 VGND.n29 VGND.t11 73.1255
R668 VGND.n32 VGND.n31 73.1255
R669 VGND.n32 VGND.t11 73.1255
R670 VGND.n144 VGND.n143 73.1255
R671 VGND.n143 VGND.t11 73.1255
R672 VGND.n147 VGND.n141 73.1255
R673 VGND.n141 VGND.t11 73.1255
R674 VGND.n124 VGND.n112 53.0829
R675 VGND.n114 VGND.n113 53.0829
R676 VGND.n118 VGND.n113 53.0829
R677 VGND.n125 VGND.n124 53.0829
R678 VGND.n133 VGND.n39 53.0829
R679 VGND.n41 VGND.n40 53.0829
R680 VGND.n45 VGND.n40 53.0829
R681 VGND.n134 VGND.n133 53.0829
R682 VGND VGND.t20 47.2522
R683 VGND.n71 VGND.t44 41.4295
R684 VGND.n71 VGND.t14 41.4295
R685 VGND.n0 VGND.t12 41.4295
R686 VGND.n0 VGND.t15 41.4295
R687 VGND.n136 VGND.t2 39.9468
R688 VGND.n128 VGND.t2 39.9468
R689 VGND.n127 VGND.t17 39.9468
R690 VGND.n119 VGND.t17 39.9468
R691 VGND.n69 VGND.n68 38.3396
R692 VGND.n19 VGND.n18 38.3396
R693 VGND.n60 VGND.n59 31.624
R694 VGND.n10 VGND.n9 31.624
R695 VGND.n65 VGND.n53 30.8711
R696 VGND.n15 VGND.n3 30.8711
R697 VGND.n61 VGND.n53 25.6005
R698 VGND.n11 VGND.n3 25.6005
R699 VGND.n52 VGND.t34 24.9236
R700 VGND.n52 VGND.t32 24.9236
R701 VGND.n55 VGND.t28 24.9236
R702 VGND.n55 VGND.t26 24.9236
R703 VGND.n66 VGND.t22 24.9236
R704 VGND.n66 VGND.t36 24.9236
R705 VGND.n2 VGND.t6 24.9236
R706 VGND.n2 VGND.t47 24.9236
R707 VGND.n5 VGND.t10 24.9236
R708 VGND.n5 VGND.t8 24.9236
R709 VGND.n16 VGND.t19 24.9236
R710 VGND.n16 VGND.t40 24.9236
R711 VGND.n61 VGND.n60 24.8476
R712 VGND.n11 VGND.n10 24.8476
R713 VGND.n67 VGND.n65 19.577
R714 VGND.n17 VGND.n15 19.577
R715 VGND.n59 VGND.n56 18.824
R716 VGND.n9 VGND.n6 18.824
R717 VGND.t16 VGND.t3 13.0569
R718 VGND.t20 VGND.t0 13.0569
R719 VGND.n95 VGND.n83 12.7179
R720 VGND.n83 VGND.n79 12.7179
R721 VGND.n92 VGND.n91 12.7179
R722 VGND.n91 VGND.n79 12.7179
R723 VGND.n88 VGND.n87 12.7179
R724 VGND.n87 VGND.n79 12.7179
R725 VGND.n85 VGND.n76 12.7179
R726 VGND.n76 VGND.n34 12.7179
R727 VGND.n101 VGND.n100 12.7179
R728 VGND.n100 VGND.n34 12.7179
R729 VGND.n84 VGND.n82 12.7179
R730 VGND.n82 VGND.n34 12.7179
R731 VGND.n152 VGND.n151 12.7179
R732 VGND.n151 VGND.n150 12.7179
R733 VGND.n142 VGND.n139 12.7179
R734 VGND.n150 VGND.n139 12.7179
R735 VGND.n149 VGND.n148 12.7179
R736 VGND.n150 VGND.n149 12.7179
R737 VGND.n155 VGND.n154 12.7179
R738 VGND.n156 VGND.n155 12.7179
R739 VGND.n158 VGND.n157 12.7179
R740 VGND.n157 VGND.n156 12.7179
R741 VGND.n146 VGND.n28 12.7179
R742 VGND.n156 VGND.n28 12.7179
R743 VGND.t3 VGND 10.8808
R744 VGND.t0 VGND 10.8808
R745 VGND.n57 VGND.n56 9.3005
R746 VGND.n59 VGND.n58 9.3005
R747 VGND.n60 VGND.n54 9.3005
R748 VGND.n62 VGND.n61 9.3005
R749 VGND.n63 VGND.n53 9.3005
R750 VGND.n65 VGND.n64 9.3005
R751 VGND.n68 VGND.n51 9.3005
R752 VGND.n7 VGND.n6 9.3005
R753 VGND.n9 VGND.n8 9.3005
R754 VGND.n10 VGND.n4 9.3005
R755 VGND.n12 VGND.n11 9.3005
R756 VGND.n13 VGND.n3 9.3005
R757 VGND.n15 VGND.n14 9.3005
R758 VGND.n18 VGND.n1 9.3005
R759 VGND.n160 VGND.n21 6.44804
R760 VGND VGND.n103 6.39894
R761 VGND.n109 VGND 4.88222
R762 VGND.n105 VGND.n104 4.54334
R763 VGND VGND.n161 3.72706
R764 VGND.n72 VGND 3.6322
R765 VGND.n70 VGND.n69 3.05653
R766 VGND.n20 VGND.n19 3.05653
R767 VGND.n104 VGND.n70 2.9055
R768 VGND.n21 VGND 2.83925
R769 VGND.n68 VGND.n67 2.25932
R770 VGND.n18 VGND.n17 2.25932
R771 VGND.n109 VGND.n21 2.08309
R772 VGND.n110 VGND.n109 2.0236
R773 VGND.n105 VGND.n38 1.8605
R774 VGND.n111 VGND.n110 1.8605
R775 VGND.n161 VGND.n160 1.85429
R776 VGND.n103 VGND.n72 1.75943
R777 VGND.n102 VGND.n101 1.35579
R778 VGND.n159 VGND.n158 1.35579
R779 VGND.n108 VGND 1.34199
R780 VGND.n107 VGND.n106 0.932201
R781 VGND.n107 VGND.n50 0.858576
R782 VGND VGND.n49 0.504285
R783 VGND VGND.n107 0.454108
R784 VGND.n72 VGND.n71 0.191676
R785 VGND.n161 VGND.n0 0.1505
R786 VGND.n64 VGND.n51 0.120292
R787 VGND.n64 VGND.n63 0.120292
R788 VGND.n63 VGND.n62 0.120292
R789 VGND.n62 VGND.n54 0.120292
R790 VGND.n58 VGND.n54 0.120292
R791 VGND.n58 VGND.n57 0.120292
R792 VGND.n14 VGND.n1 0.120292
R793 VGND.n14 VGND.n13 0.120292
R794 VGND.n13 VGND.n12 0.120292
R795 VGND.n12 VGND.n4 0.120292
R796 VGND.n8 VGND.n4 0.120292
R797 VGND.n8 VGND.n7 0.120292
R798 VGND.n20 VGND.n1 0.112479
R799 VGND.n70 VGND.n51 0.111177
R800 VGND.n106 VGND.n105 0.0971495
R801 VGND.n110 VGND.n108 0.0971495
R802 VGND.n103 VGND.n102 0.0674065
R803 VGND.n160 VGND.n159 0.0674065
R804 VGND.n57 VGND 0.0603958
R805 VGND.n7 VGND 0.0603958
R806 VGND.n50 VGND 0.0578348
R807 VGND.n49 VGND 0.0578348
R808 VGND.n104 VGND 0.0484911
R809 VGND.n20 VGND 0.0252396
R810 VGND.n70 VGND 0.0239375
R811 VGND.n70 VGND 0.02175
R812 VGND VGND.n20 0.02175
R813 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n14 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t13 212.081
R814 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n13 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t12 212.081
R815 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n1 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t11 212.081
R816 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n10 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t7 212.081
R817 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n2 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t5 212.081
R818 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n7 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t17 212.081
R819 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n5 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t16 212.081
R820 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n3 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t10 212.081
R821 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n4 tdc_0.sky130_fd_sc_hd__inv_8_1.A 171.969
R822 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n6 tdc_0.sky130_fd_sc_hd__inv_8_1.A 152
R823 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n0 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n8 152
R824 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n9 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n0 152
R825 tdc_0.sky130_fd_sc_hd__inv_8_1.A tdc_0.sky130_fd_sc_hd__inv_8_1.A.n11 152
R826 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n12 tdc_0.sky130_fd_sc_hd__inv_8_1.A 152
R827 tdc_0.sky130_fd_sc_hd__inv_8_1.A tdc_0.sky130_fd_sc_hd__inv_8_1.A.n15 152
R828 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n14 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t6 139.78
R829 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n13 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t4 139.78
R830 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n1 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t3 139.78
R831 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n10 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t15 139.78
R832 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n2 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t14 139.78
R833 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n7 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t9 139.78
R834 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n5 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t8 139.78
R835 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n3 tdc_0.sky130_fd_sc_hd__inv_8_1.A.t2 139.78
R836 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n0 tdc_0.sky130_fd_sc_hd__inv_8_1.A 44.5445
R837 tdc_0.sky130_fd_sc_hd__inv_8_1.A tdc_0.sky130_fd_sc_hd__inv_8_1.A.t0 42.5188
R838 tdc_0.sky130_fd_sc_hd__inv_8_1.A tdc_0.sky130_fd_sc_hd__inv_8_1.A.t1 39.7543
R839 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n4 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n3 30.6732
R840 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n5 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n4 30.6732
R841 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n6 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n5 30.6732
R842 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n7 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n6 30.6732
R843 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n8 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n7 30.6732
R844 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n8 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n2 30.6732
R845 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n9 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n2 30.6732
R846 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n10 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n9 30.6732
R847 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n11 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n10 30.6732
R848 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n11 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n1 30.6732
R849 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n12 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n1 30.6732
R850 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n13 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n12 30.6732
R851 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n15 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n13 30.6732
R852 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n15 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n14 30.6732
R853 tdc_0.sky130_fd_sc_hd__inv_8_1.A.n0 tdc_0.sky130_fd_sc_hd__inv_8_1.A 26.7409
R854 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n0 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t18 732.475
R855 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n0 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t17 725.527
R856 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t17 tdc_0.sky130_fd_sc_hd__inv_8_1.Y 721.894
R857 tdc_0.sky130_fd_sc_hd__inv_8_1.Y tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t16 397.69
R858 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n7 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n2 205.28
R859 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n9 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n8 205.28
R860 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n4 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n3 205.28
R861 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n6 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n5 205.28
R862 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n11 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n10 99.1749
R863 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n13 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n12 99.1749
R864 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n15 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n14 99.1749
R865 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n17 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n16 99.1749
R866 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n9 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n7 38.4005
R867 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n6 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n4 38.4005
R868 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n7 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n6 38.4005
R869 tdc_0.sky130_fd_sc_hd__inv_8_1.Y tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n9 34.4358
R870 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n13 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n11 34.3584
R871 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n15 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n13 34.3584
R872 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n17 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n15 34.3584
R873 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n4 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n1 33.2936
R874 tdc_0.sky130_fd_sc_hd__inv_8_1.Y tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n17 27.7875
R875 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n2 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t14 26.5955
R876 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n2 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t12 26.5955
R877 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n8 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t11 26.5955
R878 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n8 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t10 26.5955
R879 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n3 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t13 26.5955
R880 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n3 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t9 26.5955
R881 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n5 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t8 26.5955
R882 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n5 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t15 26.5955
R883 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n11 tdc_0.sky130_fd_sc_hd__inv_8_1.Y 25.611
R884 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n10 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t5 24.9236
R885 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n10 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t4 24.9236
R886 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n12 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t0 24.9236
R887 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n12 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t6 24.9236
R888 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n14 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t2 24.9236
R889 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n14 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t1 24.9236
R890 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n16 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t7 24.9236
R891 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n16 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t3 24.9236
R892 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n1 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n0 18.432
R893 tdc_0.sky130_fd_sc_hd__inv_8_1.Y tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n1 3.15412
R894 a_26743_17057.t0 a_26743_17057.t1 168.275
R895 ua[0] ua[0].t0 22.1303
R896 ua[0] ua[0].t1 15.5512
R897 ua[0].n0 ua[0] 14.1849
R898 ua[0].n1 ua[0] 8.94647
R899 ua[0].n1 ua[0].n0 0.906627
R900 ua[0].n0 ua[0] 0.614562
R901 ua[0] ua[0].n1 0.0311373
R902 a_25988_7882.t0 a_25988_7882.t1 80.0316
R903 a_23058_11167.t0 a_23058_11167.t1 84.355
R904 a_25891_11454.t2 a_25891_11454.t0 42.8857
R905 a_25891_11454.t1 a_25891_11454.t2 41.1012
R906 a_25891_11454.t2 a_25891_11454.t3 31.2853
R907 a_27981_11167.t0 a_27981_11167.t1 84.355
R908 a_25914_16928.t0 a_25914_16928.t1 49.8467
R909 clk.n1 clk 39.6347
R910 clk.n0 clk.t0 19.3818
R911 clk.n2 clk.t3 19.3818
R912 clk.n0 clk.t2 12.1478
R913 clk.n2 clk.t1 12.1478
R914 clk clk.n0 4.76092
R915 clk clk.n2 4.76092
R916 clk.n3 clk 4.1447
R917 clk.n3 clk.n1 2.89112
R918 clk clk.n3 2.78331
R919 clk.n1 clk 0.551542
R920 a_24477_17057.t0 a_24477_17057.t1 168.275
R921 a_26334_16003.t0 a_26334_16003.t1 169.548
R922 a_22970_11453.t3 a_22970_11453.t0 42.8857
R923 a_22970_11453.t1 a_22970_11453.t3 41.1012
R924 a_22970_11453.t3 a_22970_11453.t2 25.3663
R925 ua[1] ua[1].t1 22.1303
R926 ua[1] ua[1].t0 15.5512
R927 ua[1].n0 ua[1] 13.8786
R928 ua[1].n1 ua[1] 8.02083
R929 ua[1].n1 ua[1].n0 1.21288
R930 ua[1].n0 ua[1] 0.308313
R931 ua[1] ua[1].n1 0.0213333
R932 a_25456_16928.t0 a_25456_16928.t1 49.8467
R933 a_24251_7882.t0 a_24251_7882.t1 80.0316
R934 a_24486_16003.t0 a_24486_16003.t1 169.548
C0 tdc_0.sky130_fd_sc_hd__inv_8_0.A tdc_0.sky130_fd_sc_hd__inv_8_1.A 0.102267f
C1 uio_oe[2] uio_oe[3] 0.031023f
C2 uio_in[0] ui_in[7] 0.031023f
C3 uo_out[0] uo_out[1] 5.75124f
C4 uo_out[3] uo_out[4] 0.031023f
C5 ui_in[5] ui_in[6] 0.031023f
C6 uio_in[2] uio_in[3] 0.031023f
C7 clk VDPWR 12.3435f
C8 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A 1.56028f
C9 uio_out[6] uio_out[7] 0.031023f
C10 ui_in[2] ui_in[3] 0.031023f
C11 uio_in[5] uio_in[6] 0.031023f
C12 uio_oe[7] uio_oe[6] 0.031023f
C13 ui_in[1] ui_in[2] 0.031023f
C14 uo_out[7] uio_out[0] 0.031023f
C15 tdc_0.sky130_fd_sc_hd__inv_8_0.A VDPWR 1.25866f
C16 uo_out[0] VDPWR 0.68802f
C17 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B uo_out[1] 0.113435f
C18 ui_in[3] ui_in[4] 0.031023f
C19 uio_out[4] uio_out[5] 0.031023f
C20 tdc_0.sky130_fd_sc_hd__inv_8_1.Y tdc_0.sky130_fd_sc_hd__inv_8_0.A 0.012114f
C21 tdc_0.sky130_fd_sc_hd__inv_8_0.Y VDPWR 2.77879f
C22 uio_in[0] uio_in[1] 0.031023f
C23 uio_oe[5] uio_oe[6] 0.031023f
C24 uio_in[4] uio_in[3] 0.031023f
C25 uio_in[4] uio_in[5] 0.031023f
C26 tdc_0.sky130_fd_sc_hd__inv_8_1.Y tdc_0.sky130_fd_sc_hd__inv_8_0.Y 0.439324f
C27 uio_in[2] uio_in[1] 0.031023f
C28 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A uo_out[1] 0.404633f
C29 uio_out[6] uio_out[5] 0.031023f
C30 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B VDPWR 2.55279f
C31 uio_oe[5] uio_oe[4] 0.031023f
C32 clk ena 0.031023f
C33 uo_out[2] uo_out[1] 0.031023f
C34 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B tdc_0.sky130_fd_sc_hd__inv_8_1.Y 0.151836f
C35 ua[0] ua[1] 1.66537f
C36 uo_out[0] uio_in[7] 0.031023f
C37 uio_oe[0] uio_oe[1] 0.031023f
C38 VDPWR tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A 2.04241f
C39 uio_out[2] uio_out[1] 0.031023f
C40 uio_oe[2] uio_oe[1] 0.031023f
C41 uio_out[0] uio_out[1] 0.031023f
C42 uio_out[7] uio_oe[0] 0.031023f
C43 uio_out[4] uio_out[3] 0.031023f
C44 VDPWR ua[1] 11.5054f
C45 tdc_0.sky130_fd_sc_hd__inv_8_1.Y tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A 0.267831f
C46 uio_out[2] uio_out[3] 0.031023f
C47 tdc_0.sky130_fd_sc_hd__inv_8_0.A tdc_0.sky130_fd_sc_hd__inv_8_0.Y 1.00224f
C48 uo_out[3] uo_out[2] 0.031023f
C49 VDPWR uo_out[1] 0.345733f
C50 VDPWR tdc_0.sky130_fd_sc_hd__inv_8_1.A 1.25677f
C51 ua[0] VDPWR 11.6956f
C52 ui_in[1] ui_in[0] 0.031023f
C53 tdc_0.sky130_fd_sc_hd__inv_8_1.Y uo_out[1] 0.016955f
C54 tdc_0.sky130_fd_sc_hd__inv_8_1.Y tdc_0.sky130_fd_sc_hd__inv_8_1.A 1.01744f
C55 ui_in[5] ui_in[4] 0.031023f
C56 uio_oe[4] uio_oe[3] 0.031023f
C57 uo_out[5] uo_out[4] 0.031023f
C58 ui_in[7] ui_in[6] 0.031023f
C59 clk rst_n 0.031023f
C60 uo_out[0] tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B 0.300447f
C61 clk ua[1] 3.26149f
C62 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B tdc_0.sky130_fd_sc_hd__inv_8_0.Y 0.26039f
C63 uo_out[6] uo_out[7] 0.031023f
C64 uo_out[6] uo_out[5] 0.031023f
C65 uio_in[6] uio_in[7] 0.031023f
C66 tdc_0.sky130_fd_sc_hd__inv_8_1.Y VDPWR 2.31781f
C67 uo_out[0] tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A 0.36853f
C68 ua[0] clk 3.49067f
C69 rst_n ui_in[0] 0.031023f
C70 tdc_0.sky130_fd_sc_hd__inv_8_0.Y tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A 0.148337f
C71 ua[2] VGND 0.146962f
C72 ua[3] VGND 0.146962f
C73 ua[4] VGND 0.146962f
C74 ua[5] VGND 0.146962f
C75 ua[6] VGND 0.146962f
C76 ua[7] VGND 0.146962f
C77 ena VGND 0.070385f
C78 rst_n VGND 0.042875f
C79 ui_in[0] VGND 0.042875f
C80 ui_in[1] VGND 0.042875f
C81 ui_in[2] VGND 0.042875f
C82 ui_in[3] VGND 0.042875f
C83 ui_in[4] VGND 0.042875f
C84 ui_in[5] VGND 0.042875f
C85 ui_in[6] VGND 0.042875f
C86 ui_in[7] VGND 0.042875f
C87 uio_in[0] VGND 0.042875f
C88 uio_in[1] VGND 0.042875f
C89 uio_in[2] VGND 0.042875f
C90 uio_in[3] VGND 0.042875f
C91 uio_in[4] VGND 0.042875f
C92 uio_in[5] VGND 0.042875f
C93 uio_in[6] VGND 0.042875f
C94 uio_in[7] VGND 0.042875f
C95 uo_out[2] VGND 0.042875f
C96 uo_out[3] VGND 0.042875f
C97 uo_out[4] VGND 0.042875f
C98 uo_out[5] VGND 0.042875f
C99 uo_out[6] VGND 0.042875f
C100 uo_out[7] VGND 0.042875f
C101 uio_out[0] VGND 0.042875f
C102 uio_out[1] VGND 0.042875f
C103 uio_out[2] VGND 0.042875f
C104 uio_out[3] VGND 0.042875f
C105 uio_out[4] VGND 0.042875f
C106 uio_out[5] VGND 0.042875f
C107 uio_out[6] VGND 0.042875f
C108 uio_out[7] VGND 0.042875f
C109 uio_oe[0] VGND 0.042875f
C110 uio_oe[1] VGND 0.042875f
C111 uio_oe[2] VGND 0.042875f
C112 uio_oe[3] VGND 0.042875f
C113 uio_oe[4] VGND 0.042875f
C114 uio_oe[5] VGND 0.042875f
C115 uio_oe[6] VGND 0.042875f
C116 uio_oe[7] VGND 0.070385f
C117 ua[1] VGND 22.573984f
C118 clk VGND 44.64292f
C119 ua[0] VGND 24.011366f
C120 uo_out[1] VGND 12.907537f
C121 uo_out[0] VGND 12.838606f
C122 VDPWR VGND 0.173672p
C123 tdc_0.sky130_fd_sc_hd__inv_8_0.A VGND 2.20632f
C124 tdc_0.sky130_fd_sc_hd__inv_8_1.A VGND 2.2055f
C125 tdc_0.sky130_fd_sc_hd__inv_8_0.Y VGND 2.092111f
C126 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B VGND 1.030628f
C127 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A VGND 1.268676f
C128 tdc_0.sky130_fd_sc_hd__inv_8_1.Y VGND 2.562836f
C129 ua[1].t1 VGND 6.43383f
C130 ua[1].t0 VGND 3.19687f
C131 ua[1].n0 VGND 0.271212f
C132 ua[1].n1 VGND 0.18139f
C133 a_22970_11453.t3 VGND 6.02326f
C134 a_22970_11453.t2 VGND 1.682f
C135 a_22970_11453.t0 VGND 0.023258f
C136 a_22970_11453.t1 VGND 0.071482f
C137 clk.t2 VGND 1.91441f
C138 clk.t0 VGND 4.28996f
C139 clk.n0 VGND 1.37086f
C140 clk.n1 VGND 1.4078f
C141 clk.t3 VGND 4.28996f
C142 clk.t1 VGND 1.91441f
C143 clk.n2 VGND 1.37086f
C144 clk.n3 VGND 0.418408f
C145 a_25891_11454.t0 VGND 0.02296f
C146 a_25891_11454.t3 VGND 5.01216f
C147 a_25891_11454.t2 VGND 2.59432f
C148 a_25891_11454.t1 VGND 0.070565f
C149 ua[0].t0 VGND 6.156f
C150 ua[0].t1 VGND 3.05882f
C151 ua[0].n0 VGND 0.264584f
C152 ua[0].n1 VGND 0.346238f
C153 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t16 VGND 0.050467f
C154 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t17 VGND 0.058564f
C155 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t18 VGND 0.082833f
C156 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n0 VGND 0.837698f
C157 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n1 VGND 0.060904f
C158 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t14 VGND 0.010615f
C159 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t12 VGND 0.010615f
C160 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n2 VGND 0.023597f
C161 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t13 VGND 0.010615f
C162 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t9 VGND 0.010615f
C163 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n3 VGND 0.023597f
C164 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n4 VGND 0.066186f
C165 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t8 VGND 0.010615f
C166 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t15 VGND 0.010615f
C167 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n5 VGND 0.023597f
C168 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n6 VGND 0.061607f
C169 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n7 VGND 0.061607f
C170 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t11 VGND 0.010615f
C171 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.t10 VGND 0.010615f
C172 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n8 VGND 0.023597f
C173 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n9 VGND 0.067996f
C174 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n10 VGND 0.015714f
C175 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n11 VGND 0.049534f
C176 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n12 VGND 0.015714f
C177 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n13 VGND 0.047056f
C178 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n14 VGND 0.015714f
C179 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n15 VGND 0.047056f
C180 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n16 VGND 0.015714f
C181 tdc_0.sky130_fd_sc_hd__inv_8_1.Y.n17 VGND 0.049825f
C182 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t16 VGND 0.405879f
C183 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t17 VGND 0.265238f
C184 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t18 VGND 0.0764f
C185 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n0 VGND 0.825826f
C186 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n1 VGND 0.050107f
C187 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t12 VGND 0.013836f
C188 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t8 VGND 0.013836f
C189 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n2 VGND 0.030758f
C190 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t13 VGND 0.013836f
C191 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t11 VGND 0.013836f
C192 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n3 VGND 0.030758f
C193 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t10 VGND 0.013836f
C194 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t9 VGND 0.013836f
C195 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n4 VGND 0.030758f
C196 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n5 VGND 0.020483f
C197 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n6 VGND 0.020483f
C198 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n7 VGND 0.020483f
C199 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n8 VGND 0.020483f
C200 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n9 VGND 0.067676f
C201 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n10 VGND 0.061337f
C202 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n11 VGND 0.061337f
C203 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n12 VGND 0.070017f
C204 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n13 VGND 0.083443f
C205 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n14 VGND 0.080303f
C206 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t7 VGND 0.013836f
C207 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.t14 VGND 0.013836f
C208 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n15 VGND 0.030757f
C209 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n16 VGND 0.080303f
C210 tdc_0.sky130_fd_sc_hd__inv_8_0.Y.n17 VGND 0.083713f
C211 uo_out[1].t4 VGND 0.011512f
C212 uo_out[1].n0 VGND 0.022651f
C213 uo_out[1].t1 VGND 0.013802f
C214 uo_out[1].n2 VGND 0.018341f
C215 uo_out[1].n4 VGND 0.012268f
C216 uo_out[1].n5 VGND 0.02452f
C217 uo_out[1].n6 VGND 0.071864f
C218 uo_out[1].n7 VGND 2.21232f
C219 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n0 VGND 1.05323f
C220 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t6 VGND 0.015592f
C221 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t3 VGND 0.024984f
C222 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n1 VGND 0.049158f
C223 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t4 VGND 0.063098f
C224 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t5 VGND 0.112699f
C225 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n2 VGND 0.3435f
C226 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t0 VGND 0.057939f
C227 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t1 VGND 0.181196f
C228 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n3 VGND 0.423038f
C229 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.t2 VGND 0.242161f
C230 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_0.B.n4 VGND 0.026911f
C231 VDPWR.n0 VGND 0.459508f
C232 VDPWR.n1 VGND 0.129808f
C233 VDPWR.n2 VGND 0.516796f
C234 VDPWR.n3 VGND 0.144179f
C235 VDPWR.n4 VGND 0.062397f
C236 VDPWR.n5 VGND 0.029069f
C237 VDPWR.n6 VGND 0.077304f
C238 VDPWR.n7 VGND 0.074092f
C239 VDPWR.n8 VGND 0.077304f
C240 VDPWR.n9 VGND 4.86954f
C241 VDPWR.n10 VGND 4.90327f
C242 VDPWR.n11 VGND 0.077747f
C243 VDPWR.n12 VGND 0.029395f
C244 VDPWR.n13 VGND 0.029395f
C245 VDPWR.n14 VGND 0.077747f
C246 VDPWR.n15 VGND 0.077304f
C247 VDPWR.n16 VGND 0.077304f
C248 VDPWR.n17 VGND 0.178435f
C249 VDPWR.n18 VGND 0.077304f
C250 VDPWR.n19 VGND 0.077747f
C251 VDPWR.t34 VGND 0.072177f
C252 VDPWR.t36 VGND 0.072177f
C253 VDPWR.n20 VGND 0.414028f
C254 VDPWR.n21 VGND 0.077747f
C255 VDPWR.n22 VGND 0.077747f
C256 VDPWR.n23 VGND 4.90327f
C257 VDPWR.n24 VGND 0.074092f
C258 VDPWR.n25 VGND 0.077304f
C259 VDPWR.n26 VGND 0.092679f
C260 VDPWR.n27 VGND 0.029395f
C261 VDPWR.t5 VGND 0.554361f
C262 VDPWR.n29 VGND 0.014853f
C263 VDPWR.n30 VGND 0.023596f
C264 VDPWR.n31 VGND 0.015005f
C265 VDPWR.n32 VGND 0.023596f
C266 VDPWR.n33 VGND 0.017883f
C267 VDPWR.n34 VGND 0.014853f
C268 VDPWR.n35 VGND 0.015005f
C269 VDPWR.n36 VGND 0.015005f
C270 VDPWR.n37 VGND 0.023596f
C271 VDPWR.t17 VGND 0.036763f
C272 VDPWR.t11 VGND 0.011604f
C273 VDPWR.t33 VGND 0.011604f
C274 VDPWR.n39 VGND 0.012461f
C275 VDPWR.n42 VGND 0.013568f
C276 VDPWR.n47 VGND 0.015334f
C277 VDPWR.t29 VGND 0.011602f
C278 VDPWR.t31 VGND 0.011602f
C279 VDPWR.n49 VGND 0.024129f
C280 VDPWR.n51 VGND 0.012461f
C281 VDPWR.n52 VGND 0.012461f
C282 VDPWR.n53 VGND 0.012461f
C283 VDPWR.n55 VGND 0.015334f
C284 VDPWR.n57 VGND 0.012461f
C285 VDPWR.n58 VGND 0.012461f
C286 VDPWR.n59 VGND 0.011309f
C287 VDPWR.n61 VGND 0.022981f
C288 VDPWR.n62 VGND 0.019546f
C289 VDPWR.t20 VGND 0.040171f
C290 VDPWR.t8 VGND 0.012154f
C291 VDPWR.n65 VGND 0.015633f
C292 VDPWR.t19 VGND 0.012158f
C293 VDPWR.n68 VGND 0.016735f
C294 VDPWR.n70 VGND 0.012362f
C295 VDPWR.t6 VGND 0.0402f
C296 VDPWR.t24 VGND 0.012154f
C297 VDPWR.n73 VGND 0.015633f
C298 VDPWR.t1 VGND 0.012158f
C299 VDPWR.n75 VGND 0.016735f
C300 VDPWR.n78 VGND 0.082582f
C301 VDPWR.n79 VGND 0.016101f
C302 VDPWR.n80 VGND 0.016071f
C303 VDPWR.n81 VGND 0.081702f
C304 VDPWR.n82 VGND 0.027089f
C305 VDPWR.t26 VGND 0.036763f
C306 VDPWR.n83 VGND 0.014853f
C307 VDPWR.n84 VGND 0.014853f
C308 VDPWR.n85 VGND 0.014853f
C309 VDPWR.n86 VGND 0.014853f
C310 VDPWR.n87 VGND 0.34023f
C311 VDPWR.t18 VGND 0.0916f
C312 VDPWR.t7 VGND 0.160003f
C313 VDPWR.n88 VGND 0.38722f
C314 VDPWR.n89 VGND 0.017883f
C315 VDPWR.n90 VGND 0.017883f
C316 VDPWR.n91 VGND 0.014853f
C317 VDPWR.n92 VGND 0.014853f
C318 VDPWR.n93 VGND 0.014853f
C319 VDPWR.n94 VGND 0.015005f
C320 VDPWR.n95 VGND 0.015005f
C321 VDPWR.n98 VGND 0.015005f
C322 VDPWR.n99 VGND 0.017883f
C323 VDPWR.n100 VGND 0.015005f
C324 VDPWR.n101 VGND 0.015005f
C325 VDPWR.n102 VGND 0.015005f
C326 VDPWR.n105 VGND 0.015005f
C327 VDPWR.n106 VGND 0.017883f
C328 VDPWR.n107 VGND 0.015005f
C329 VDPWR.n108 VGND 0.014853f
C330 VDPWR.n109 VGND 0.023596f
C331 VDPWR.n110 VGND 0.023596f
C332 VDPWR.t4 VGND 0.554361f
C333 VDPWR.n111 VGND 0.023596f
C334 VDPWR.n112 VGND 0.044825f
C335 VDPWR.n113 VGND 0.142536f
C336 VDPWR.n114 VGND 0.054602f
C337 VDPWR.n115 VGND 0.058131f
C338 VDPWR.n116 VGND 0.158083f
C339 VDPWR.n117 VGND 0.044825f
C340 VDPWR.n118 VGND 0.014853f
C341 VDPWR.n119 VGND 0.014853f
C342 VDPWR.n120 VGND 0.017883f
C343 VDPWR.n121 VGND 0.015005f
C344 VDPWR.n123 VGND 0.015005f
C345 VDPWR.n124 VGND 0.014853f
C346 VDPWR.n125 VGND 0.014853f
C347 VDPWR.n126 VGND 0.34023f
C348 VDPWR.n128 VGND 0.015005f
C349 VDPWR.n129 VGND 0.017883f
C350 VDPWR.n130 VGND 0.017883f
C351 VDPWR.n131 VGND 0.015005f
C352 VDPWR.n133 VGND 0.015005f
C353 VDPWR.n134 VGND 0.014853f
C354 VDPWR.n135 VGND 0.014853f
C355 VDPWR.n136 VGND 0.347963f
C356 VDPWR.t0 VGND 0.0916f
C357 VDPWR.t23 VGND 0.163734f
C358 VDPWR.t9 VGND 0.266485f
C359 VDPWR.t13 VGND 0.255674f
C360 VDPWR.n137 VGND 1.42639f
C361 VDPWR.n138 VGND 4.89765f
C362 VDPWR.n139 VGND 0.077304f
C363 VDPWR.n140 VGND 0.062397f
C364 VDPWR.n141 VGND 0.077747f
C365 VDPWR.n142 VGND 0.077304f
C366 VDPWR.n143 VGND 0.074092f
C367 VDPWR.n144 VGND 0.077747f
C368 VDPWR.n145 VGND 0.062397f
C369 VDPWR.n146 VGND 0.062397f
C370 VDPWR.n147 VGND 0.077747f
C371 VDPWR.n148 VGND 0.029069f
C372 VDPWR.n149 VGND 0.144179f
C373 VDPWR.n150 VGND 0.160967f
C374 VDPWR.n151 VGND 0.178476f
C375 VDPWR.n152 VGND 0.092679f
C376 VDPWR.t21 VGND 8.61447f
C377 VDPWR.n153 VGND 0.029395f
C378 VDPWR.n154 VGND 0.029069f
C379 VDPWR.n155 VGND 0.144179f
C380 VDPWR.n156 VGND 0.161007f
C381 VDPWR.n157 VGND 0.360761f
C382 VDPWR.n158 VGND 0.161007f
C383 VDPWR.n159 VGND 0.077747f
C384 VDPWR.n160 VGND 0.077747f
C385 VDPWR.n161 VGND 0.077747f
C386 VDPWR.n162 VGND 0.062397f
C387 VDPWR.n163 VGND 0.062397f
C388 VDPWR.t28 VGND 0.072177f
C389 VDPWR.t3 VGND 0.072177f
C390 VDPWR.n164 VGND 0.414028f
C391 VDPWR.n165 VGND 0.029069f
C392 VDPWR.n166 VGND 0.077747f
C393 VDPWR.n167 VGND 0.074092f
C394 VDPWR.n168 VGND 0.178435f
C395 VDPWR.n169 VGND 0.092679f
C396 VDPWR.t2 VGND 8.61447f
C397 VDPWR.n170 VGND 0.092679f
C398 VDPWR.n171 VGND 0.178435f
C399 VDPWR.n172 VGND 0.161007f
C400 VDPWR.n173 VGND 0.144179f
C401 VDPWR.n174 VGND 0.129808f
C402 VDPWR.n175 VGND 0.397175f
C403 VDPWR.n176 VGND 1.2257f
C404 uo_out[0].t1 VGND 0.013561f
C405 uo_out[0].n0 VGND 0.0139f
C406 uo_out[0].t4 VGND 0.011325f
C407 uo_out[0].n1 VGND 0.021557f
C408 uo_out[0].n2 VGND 0.064611f
C409 uo_out[0].n3 VGND 0.06413f
C410 uo_out[0].n5 VGND 0.012053f
C411 uo_out[0].n6 VGND 0.02863f
C412 uo_out[0].n7 VGND 2.21241f
C413 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n0 VGND 0.822986f
C414 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t6 VGND 0.01191f
C415 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t3 VGND 0.019075f
C416 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n1 VGND 0.036309f
C417 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t0 VGND 0.043796f
C418 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t2 VGND 0.138855f
C419 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n2 VGND 0.322247f
C420 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t1 VGND 0.186869f
C421 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t4 VGND 0.048052f
C422 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.t5 VGND 0.085969f
C423 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n3 VGND 0.261649f
C424 tdc_0.phase_detector_0.sky130_fd_sc_hd__nand2_1_1.A.n4 VGND 0.016138f
.ends

