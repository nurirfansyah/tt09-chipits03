magic
tech sky130A
magscale 1 2
timestamp 1729057844
<< error_p >>
rect -29 572 29 578
rect -29 538 -17 572
rect -29 532 29 538
rect -29 -538 29 -532
rect -29 -572 -17 -538
rect -29 -578 29 -572
<< pwell >>
rect -226 -710 226 710
<< nmos >>
rect -30 -500 30 500
<< ndiff >>
rect -88 488 -30 500
rect -88 -488 -76 488
rect -42 -488 -30 488
rect -88 -500 -30 -488
rect 30 488 88 500
rect 30 -488 42 488
rect 76 -488 88 488
rect 30 -500 88 -488
<< ndiffc >>
rect -76 -488 -42 488
rect 42 -488 76 488
<< psubdiff >>
rect -190 640 -94 674
rect 94 640 190 674
rect -190 578 -156 640
rect 156 578 190 640
rect -190 -640 -156 -578
rect 156 -640 190 -578
rect -190 -674 -94 -640
rect 94 -674 190 -640
<< psubdiffcont >>
rect -94 640 94 674
rect -190 -578 -156 578
rect 156 -578 190 578
rect -94 -674 94 -640
<< poly >>
rect -33 572 33 588
rect -33 538 -17 572
rect 17 538 33 572
rect -33 522 33 538
rect -30 500 30 522
rect -30 -522 30 -500
rect -33 -538 33 -522
rect -33 -572 -17 -538
rect 17 -572 33 -538
rect -33 -588 33 -572
<< polycont >>
rect -17 538 17 572
rect -17 -572 17 -538
<< locali >>
rect -190 640 -94 674
rect 94 640 190 674
rect -190 578 -156 640
rect 156 578 190 640
rect -33 538 -17 572
rect 17 538 33 572
rect -76 488 -42 504
rect -76 -504 -42 -488
rect 42 488 76 504
rect 42 -504 76 -488
rect -33 -572 -17 -538
rect 17 -572 33 -538
rect -190 -640 -156 -578
rect 156 -640 190 -578
rect -190 -674 -94 -640
rect 94 -674 190 -640
<< viali >>
rect -17 538 17 572
rect -76 -488 -42 488
rect 42 -488 76 488
rect -17 -572 17 -538
<< metal1 >>
rect -29 572 29 578
rect -29 538 -17 572
rect 17 538 29 572
rect -29 532 29 538
rect -82 488 -36 500
rect -82 -488 -76 488
rect -42 -488 -36 488
rect -82 -500 -36 -488
rect 36 488 82 500
rect 36 -488 42 488
rect 76 -488 82 488
rect 36 -500 82 -488
rect -29 -538 29 -532
rect -29 -572 -17 -538
rect 17 -572 29 -538
rect -29 -578 29 -572
<< properties >>
string FIXED_BBOX -173 -657 173 657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
