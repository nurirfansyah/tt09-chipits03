magic
tech sky130A
magscale 1 2
timestamp 1730269323
<< metal3 >>
rect -386 22892 386 22920
rect -386 22468 302 22892
rect 366 22468 386 22892
rect -386 22440 386 22468
rect -386 22172 386 22200
rect -386 21748 302 22172
rect 366 21748 386 22172
rect -386 21720 386 21748
rect -386 21452 386 21480
rect -386 21028 302 21452
rect 366 21028 386 21452
rect -386 21000 386 21028
rect -386 20732 386 20760
rect -386 20308 302 20732
rect 366 20308 386 20732
rect -386 20280 386 20308
rect -386 20012 386 20040
rect -386 19588 302 20012
rect 366 19588 386 20012
rect -386 19560 386 19588
rect -386 19292 386 19320
rect -386 18868 302 19292
rect 366 18868 386 19292
rect -386 18840 386 18868
rect -386 18572 386 18600
rect -386 18148 302 18572
rect 366 18148 386 18572
rect -386 18120 386 18148
rect -386 17852 386 17880
rect -386 17428 302 17852
rect 366 17428 386 17852
rect -386 17400 386 17428
rect -386 17132 386 17160
rect -386 16708 302 17132
rect 366 16708 386 17132
rect -386 16680 386 16708
rect -386 16412 386 16440
rect -386 15988 302 16412
rect 366 15988 386 16412
rect -386 15960 386 15988
rect -386 15692 386 15720
rect -386 15268 302 15692
rect 366 15268 386 15692
rect -386 15240 386 15268
rect -386 14972 386 15000
rect -386 14548 302 14972
rect 366 14548 386 14972
rect -386 14520 386 14548
rect -386 14252 386 14280
rect -386 13828 302 14252
rect 366 13828 386 14252
rect -386 13800 386 13828
rect -386 13532 386 13560
rect -386 13108 302 13532
rect 366 13108 386 13532
rect -386 13080 386 13108
rect -386 12812 386 12840
rect -386 12388 302 12812
rect 366 12388 386 12812
rect -386 12360 386 12388
rect -386 12092 386 12120
rect -386 11668 302 12092
rect 366 11668 386 12092
rect -386 11640 386 11668
rect -386 11372 386 11400
rect -386 10948 302 11372
rect 366 10948 386 11372
rect -386 10920 386 10948
rect -386 10652 386 10680
rect -386 10228 302 10652
rect 366 10228 386 10652
rect -386 10200 386 10228
rect -386 9932 386 9960
rect -386 9508 302 9932
rect 366 9508 386 9932
rect -386 9480 386 9508
rect -386 9212 386 9240
rect -386 8788 302 9212
rect 366 8788 386 9212
rect -386 8760 386 8788
rect -386 8492 386 8520
rect -386 8068 302 8492
rect 366 8068 386 8492
rect -386 8040 386 8068
rect -386 7772 386 7800
rect -386 7348 302 7772
rect 366 7348 386 7772
rect -386 7320 386 7348
rect -386 7052 386 7080
rect -386 6628 302 7052
rect 366 6628 386 7052
rect -386 6600 386 6628
rect -386 6332 386 6360
rect -386 5908 302 6332
rect 366 5908 386 6332
rect -386 5880 386 5908
rect -386 5612 386 5640
rect -386 5188 302 5612
rect 366 5188 386 5612
rect -386 5160 386 5188
rect -386 4892 386 4920
rect -386 4468 302 4892
rect 366 4468 386 4892
rect -386 4440 386 4468
rect -386 4172 386 4200
rect -386 3748 302 4172
rect 366 3748 386 4172
rect -386 3720 386 3748
rect -386 3452 386 3480
rect -386 3028 302 3452
rect 366 3028 386 3452
rect -386 3000 386 3028
rect -386 2732 386 2760
rect -386 2308 302 2732
rect 366 2308 386 2732
rect -386 2280 386 2308
rect -386 2012 386 2040
rect -386 1588 302 2012
rect 366 1588 386 2012
rect -386 1560 386 1588
rect -386 1292 386 1320
rect -386 868 302 1292
rect 366 868 386 1292
rect -386 840 386 868
rect -386 572 386 600
rect -386 148 302 572
rect 366 148 386 572
rect -386 120 386 148
rect -386 -148 386 -120
rect -386 -572 302 -148
rect 366 -572 386 -148
rect -386 -600 386 -572
rect -386 -868 386 -840
rect -386 -1292 302 -868
rect 366 -1292 386 -868
rect -386 -1320 386 -1292
rect -386 -1588 386 -1560
rect -386 -2012 302 -1588
rect 366 -2012 386 -1588
rect -386 -2040 386 -2012
rect -386 -2308 386 -2280
rect -386 -2732 302 -2308
rect 366 -2732 386 -2308
rect -386 -2760 386 -2732
rect -386 -3028 386 -3000
rect -386 -3452 302 -3028
rect 366 -3452 386 -3028
rect -386 -3480 386 -3452
rect -386 -3748 386 -3720
rect -386 -4172 302 -3748
rect 366 -4172 386 -3748
rect -386 -4200 386 -4172
rect -386 -4468 386 -4440
rect -386 -4892 302 -4468
rect 366 -4892 386 -4468
rect -386 -4920 386 -4892
rect -386 -5188 386 -5160
rect -386 -5612 302 -5188
rect 366 -5612 386 -5188
rect -386 -5640 386 -5612
rect -386 -5908 386 -5880
rect -386 -6332 302 -5908
rect 366 -6332 386 -5908
rect -386 -6360 386 -6332
rect -386 -6628 386 -6600
rect -386 -7052 302 -6628
rect 366 -7052 386 -6628
rect -386 -7080 386 -7052
rect -386 -7348 386 -7320
rect -386 -7772 302 -7348
rect 366 -7772 386 -7348
rect -386 -7800 386 -7772
rect -386 -8068 386 -8040
rect -386 -8492 302 -8068
rect 366 -8492 386 -8068
rect -386 -8520 386 -8492
rect -386 -8788 386 -8760
rect -386 -9212 302 -8788
rect 366 -9212 386 -8788
rect -386 -9240 386 -9212
rect -386 -9508 386 -9480
rect -386 -9932 302 -9508
rect 366 -9932 386 -9508
rect -386 -9960 386 -9932
rect -386 -10228 386 -10200
rect -386 -10652 302 -10228
rect 366 -10652 386 -10228
rect -386 -10680 386 -10652
rect -386 -10948 386 -10920
rect -386 -11372 302 -10948
rect 366 -11372 386 -10948
rect -386 -11400 386 -11372
rect -386 -11668 386 -11640
rect -386 -12092 302 -11668
rect 366 -12092 386 -11668
rect -386 -12120 386 -12092
rect -386 -12388 386 -12360
rect -386 -12812 302 -12388
rect 366 -12812 386 -12388
rect -386 -12840 386 -12812
rect -386 -13108 386 -13080
rect -386 -13532 302 -13108
rect 366 -13532 386 -13108
rect -386 -13560 386 -13532
rect -386 -13828 386 -13800
rect -386 -14252 302 -13828
rect 366 -14252 386 -13828
rect -386 -14280 386 -14252
rect -386 -14548 386 -14520
rect -386 -14972 302 -14548
rect 366 -14972 386 -14548
rect -386 -15000 386 -14972
rect -386 -15268 386 -15240
rect -386 -15692 302 -15268
rect 366 -15692 386 -15268
rect -386 -15720 386 -15692
rect -386 -15988 386 -15960
rect -386 -16412 302 -15988
rect 366 -16412 386 -15988
rect -386 -16440 386 -16412
rect -386 -16708 386 -16680
rect -386 -17132 302 -16708
rect 366 -17132 386 -16708
rect -386 -17160 386 -17132
rect -386 -17428 386 -17400
rect -386 -17852 302 -17428
rect 366 -17852 386 -17428
rect -386 -17880 386 -17852
rect -386 -18148 386 -18120
rect -386 -18572 302 -18148
rect 366 -18572 386 -18148
rect -386 -18600 386 -18572
rect -386 -18868 386 -18840
rect -386 -19292 302 -18868
rect 366 -19292 386 -18868
rect -386 -19320 386 -19292
rect -386 -19588 386 -19560
rect -386 -20012 302 -19588
rect 366 -20012 386 -19588
rect -386 -20040 386 -20012
rect -386 -20308 386 -20280
rect -386 -20732 302 -20308
rect 366 -20732 386 -20308
rect -386 -20760 386 -20732
rect -386 -21028 386 -21000
rect -386 -21452 302 -21028
rect 366 -21452 386 -21028
rect -386 -21480 386 -21452
rect -386 -21748 386 -21720
rect -386 -22172 302 -21748
rect 366 -22172 386 -21748
rect -386 -22200 386 -22172
rect -386 -22468 386 -22440
rect -386 -22892 302 -22468
rect 366 -22892 386 -22468
rect -386 -22920 386 -22892
<< via3 >>
rect 302 22468 366 22892
rect 302 21748 366 22172
rect 302 21028 366 21452
rect 302 20308 366 20732
rect 302 19588 366 20012
rect 302 18868 366 19292
rect 302 18148 366 18572
rect 302 17428 366 17852
rect 302 16708 366 17132
rect 302 15988 366 16412
rect 302 15268 366 15692
rect 302 14548 366 14972
rect 302 13828 366 14252
rect 302 13108 366 13532
rect 302 12388 366 12812
rect 302 11668 366 12092
rect 302 10948 366 11372
rect 302 10228 366 10652
rect 302 9508 366 9932
rect 302 8788 366 9212
rect 302 8068 366 8492
rect 302 7348 366 7772
rect 302 6628 366 7052
rect 302 5908 366 6332
rect 302 5188 366 5612
rect 302 4468 366 4892
rect 302 3748 366 4172
rect 302 3028 366 3452
rect 302 2308 366 2732
rect 302 1588 366 2012
rect 302 868 366 1292
rect 302 148 366 572
rect 302 -572 366 -148
rect 302 -1292 366 -868
rect 302 -2012 366 -1588
rect 302 -2732 366 -2308
rect 302 -3452 366 -3028
rect 302 -4172 366 -3748
rect 302 -4892 366 -4468
rect 302 -5612 366 -5188
rect 302 -6332 366 -5908
rect 302 -7052 366 -6628
rect 302 -7772 366 -7348
rect 302 -8492 366 -8068
rect 302 -9212 366 -8788
rect 302 -9932 366 -9508
rect 302 -10652 366 -10228
rect 302 -11372 366 -10948
rect 302 -12092 366 -11668
rect 302 -12812 366 -12388
rect 302 -13532 366 -13108
rect 302 -14252 366 -13828
rect 302 -14972 366 -14548
rect 302 -15692 366 -15268
rect 302 -16412 366 -15988
rect 302 -17132 366 -16708
rect 302 -17852 366 -17428
rect 302 -18572 366 -18148
rect 302 -19292 366 -18868
rect 302 -20012 366 -19588
rect 302 -20732 366 -20308
rect 302 -21452 366 -21028
rect 302 -22172 366 -21748
rect 302 -22892 366 -22468
<< mimcap >>
rect -346 22840 54 22880
rect -346 22520 -306 22840
rect 14 22520 54 22840
rect -346 22480 54 22520
rect -346 22120 54 22160
rect -346 21800 -306 22120
rect 14 21800 54 22120
rect -346 21760 54 21800
rect -346 21400 54 21440
rect -346 21080 -306 21400
rect 14 21080 54 21400
rect -346 21040 54 21080
rect -346 20680 54 20720
rect -346 20360 -306 20680
rect 14 20360 54 20680
rect -346 20320 54 20360
rect -346 19960 54 20000
rect -346 19640 -306 19960
rect 14 19640 54 19960
rect -346 19600 54 19640
rect -346 19240 54 19280
rect -346 18920 -306 19240
rect 14 18920 54 19240
rect -346 18880 54 18920
rect -346 18520 54 18560
rect -346 18200 -306 18520
rect 14 18200 54 18520
rect -346 18160 54 18200
rect -346 17800 54 17840
rect -346 17480 -306 17800
rect 14 17480 54 17800
rect -346 17440 54 17480
rect -346 17080 54 17120
rect -346 16760 -306 17080
rect 14 16760 54 17080
rect -346 16720 54 16760
rect -346 16360 54 16400
rect -346 16040 -306 16360
rect 14 16040 54 16360
rect -346 16000 54 16040
rect -346 15640 54 15680
rect -346 15320 -306 15640
rect 14 15320 54 15640
rect -346 15280 54 15320
rect -346 14920 54 14960
rect -346 14600 -306 14920
rect 14 14600 54 14920
rect -346 14560 54 14600
rect -346 14200 54 14240
rect -346 13880 -306 14200
rect 14 13880 54 14200
rect -346 13840 54 13880
rect -346 13480 54 13520
rect -346 13160 -306 13480
rect 14 13160 54 13480
rect -346 13120 54 13160
rect -346 12760 54 12800
rect -346 12440 -306 12760
rect 14 12440 54 12760
rect -346 12400 54 12440
rect -346 12040 54 12080
rect -346 11720 -306 12040
rect 14 11720 54 12040
rect -346 11680 54 11720
rect -346 11320 54 11360
rect -346 11000 -306 11320
rect 14 11000 54 11320
rect -346 10960 54 11000
rect -346 10600 54 10640
rect -346 10280 -306 10600
rect 14 10280 54 10600
rect -346 10240 54 10280
rect -346 9880 54 9920
rect -346 9560 -306 9880
rect 14 9560 54 9880
rect -346 9520 54 9560
rect -346 9160 54 9200
rect -346 8840 -306 9160
rect 14 8840 54 9160
rect -346 8800 54 8840
rect -346 8440 54 8480
rect -346 8120 -306 8440
rect 14 8120 54 8440
rect -346 8080 54 8120
rect -346 7720 54 7760
rect -346 7400 -306 7720
rect 14 7400 54 7720
rect -346 7360 54 7400
rect -346 7000 54 7040
rect -346 6680 -306 7000
rect 14 6680 54 7000
rect -346 6640 54 6680
rect -346 6280 54 6320
rect -346 5960 -306 6280
rect 14 5960 54 6280
rect -346 5920 54 5960
rect -346 5560 54 5600
rect -346 5240 -306 5560
rect 14 5240 54 5560
rect -346 5200 54 5240
rect -346 4840 54 4880
rect -346 4520 -306 4840
rect 14 4520 54 4840
rect -346 4480 54 4520
rect -346 4120 54 4160
rect -346 3800 -306 4120
rect 14 3800 54 4120
rect -346 3760 54 3800
rect -346 3400 54 3440
rect -346 3080 -306 3400
rect 14 3080 54 3400
rect -346 3040 54 3080
rect -346 2680 54 2720
rect -346 2360 -306 2680
rect 14 2360 54 2680
rect -346 2320 54 2360
rect -346 1960 54 2000
rect -346 1640 -306 1960
rect 14 1640 54 1960
rect -346 1600 54 1640
rect -346 1240 54 1280
rect -346 920 -306 1240
rect 14 920 54 1240
rect -346 880 54 920
rect -346 520 54 560
rect -346 200 -306 520
rect 14 200 54 520
rect -346 160 54 200
rect -346 -200 54 -160
rect -346 -520 -306 -200
rect 14 -520 54 -200
rect -346 -560 54 -520
rect -346 -920 54 -880
rect -346 -1240 -306 -920
rect 14 -1240 54 -920
rect -346 -1280 54 -1240
rect -346 -1640 54 -1600
rect -346 -1960 -306 -1640
rect 14 -1960 54 -1640
rect -346 -2000 54 -1960
rect -346 -2360 54 -2320
rect -346 -2680 -306 -2360
rect 14 -2680 54 -2360
rect -346 -2720 54 -2680
rect -346 -3080 54 -3040
rect -346 -3400 -306 -3080
rect 14 -3400 54 -3080
rect -346 -3440 54 -3400
rect -346 -3800 54 -3760
rect -346 -4120 -306 -3800
rect 14 -4120 54 -3800
rect -346 -4160 54 -4120
rect -346 -4520 54 -4480
rect -346 -4840 -306 -4520
rect 14 -4840 54 -4520
rect -346 -4880 54 -4840
rect -346 -5240 54 -5200
rect -346 -5560 -306 -5240
rect 14 -5560 54 -5240
rect -346 -5600 54 -5560
rect -346 -5960 54 -5920
rect -346 -6280 -306 -5960
rect 14 -6280 54 -5960
rect -346 -6320 54 -6280
rect -346 -6680 54 -6640
rect -346 -7000 -306 -6680
rect 14 -7000 54 -6680
rect -346 -7040 54 -7000
rect -346 -7400 54 -7360
rect -346 -7720 -306 -7400
rect 14 -7720 54 -7400
rect -346 -7760 54 -7720
rect -346 -8120 54 -8080
rect -346 -8440 -306 -8120
rect 14 -8440 54 -8120
rect -346 -8480 54 -8440
rect -346 -8840 54 -8800
rect -346 -9160 -306 -8840
rect 14 -9160 54 -8840
rect -346 -9200 54 -9160
rect -346 -9560 54 -9520
rect -346 -9880 -306 -9560
rect 14 -9880 54 -9560
rect -346 -9920 54 -9880
rect -346 -10280 54 -10240
rect -346 -10600 -306 -10280
rect 14 -10600 54 -10280
rect -346 -10640 54 -10600
rect -346 -11000 54 -10960
rect -346 -11320 -306 -11000
rect 14 -11320 54 -11000
rect -346 -11360 54 -11320
rect -346 -11720 54 -11680
rect -346 -12040 -306 -11720
rect 14 -12040 54 -11720
rect -346 -12080 54 -12040
rect -346 -12440 54 -12400
rect -346 -12760 -306 -12440
rect 14 -12760 54 -12440
rect -346 -12800 54 -12760
rect -346 -13160 54 -13120
rect -346 -13480 -306 -13160
rect 14 -13480 54 -13160
rect -346 -13520 54 -13480
rect -346 -13880 54 -13840
rect -346 -14200 -306 -13880
rect 14 -14200 54 -13880
rect -346 -14240 54 -14200
rect -346 -14600 54 -14560
rect -346 -14920 -306 -14600
rect 14 -14920 54 -14600
rect -346 -14960 54 -14920
rect -346 -15320 54 -15280
rect -346 -15640 -306 -15320
rect 14 -15640 54 -15320
rect -346 -15680 54 -15640
rect -346 -16040 54 -16000
rect -346 -16360 -306 -16040
rect 14 -16360 54 -16040
rect -346 -16400 54 -16360
rect -346 -16760 54 -16720
rect -346 -17080 -306 -16760
rect 14 -17080 54 -16760
rect -346 -17120 54 -17080
rect -346 -17480 54 -17440
rect -346 -17800 -306 -17480
rect 14 -17800 54 -17480
rect -346 -17840 54 -17800
rect -346 -18200 54 -18160
rect -346 -18520 -306 -18200
rect 14 -18520 54 -18200
rect -346 -18560 54 -18520
rect -346 -18920 54 -18880
rect -346 -19240 -306 -18920
rect 14 -19240 54 -18920
rect -346 -19280 54 -19240
rect -346 -19640 54 -19600
rect -346 -19960 -306 -19640
rect 14 -19960 54 -19640
rect -346 -20000 54 -19960
rect -346 -20360 54 -20320
rect -346 -20680 -306 -20360
rect 14 -20680 54 -20360
rect -346 -20720 54 -20680
rect -346 -21080 54 -21040
rect -346 -21400 -306 -21080
rect 14 -21400 54 -21080
rect -346 -21440 54 -21400
rect -346 -21800 54 -21760
rect -346 -22120 -306 -21800
rect 14 -22120 54 -21800
rect -346 -22160 54 -22120
rect -346 -22520 54 -22480
rect -346 -22840 -306 -22520
rect 14 -22840 54 -22520
rect -346 -22880 54 -22840
<< mimcapcontact >>
rect -306 22520 14 22840
rect -306 21800 14 22120
rect -306 21080 14 21400
rect -306 20360 14 20680
rect -306 19640 14 19960
rect -306 18920 14 19240
rect -306 18200 14 18520
rect -306 17480 14 17800
rect -306 16760 14 17080
rect -306 16040 14 16360
rect -306 15320 14 15640
rect -306 14600 14 14920
rect -306 13880 14 14200
rect -306 13160 14 13480
rect -306 12440 14 12760
rect -306 11720 14 12040
rect -306 11000 14 11320
rect -306 10280 14 10600
rect -306 9560 14 9880
rect -306 8840 14 9160
rect -306 8120 14 8440
rect -306 7400 14 7720
rect -306 6680 14 7000
rect -306 5960 14 6280
rect -306 5240 14 5560
rect -306 4520 14 4840
rect -306 3800 14 4120
rect -306 3080 14 3400
rect -306 2360 14 2680
rect -306 1640 14 1960
rect -306 920 14 1240
rect -306 200 14 520
rect -306 -520 14 -200
rect -306 -1240 14 -920
rect -306 -1960 14 -1640
rect -306 -2680 14 -2360
rect -306 -3400 14 -3080
rect -306 -4120 14 -3800
rect -306 -4840 14 -4520
rect -306 -5560 14 -5240
rect -306 -6280 14 -5960
rect -306 -7000 14 -6680
rect -306 -7720 14 -7400
rect -306 -8440 14 -8120
rect -306 -9160 14 -8840
rect -306 -9880 14 -9560
rect -306 -10600 14 -10280
rect -306 -11320 14 -11000
rect -306 -12040 14 -11720
rect -306 -12760 14 -12440
rect -306 -13480 14 -13160
rect -306 -14200 14 -13880
rect -306 -14920 14 -14600
rect -306 -15640 14 -15320
rect -306 -16360 14 -16040
rect -306 -17080 14 -16760
rect -306 -17800 14 -17480
rect -306 -18520 14 -18200
rect -306 -19240 14 -18920
rect -306 -19960 14 -19640
rect -306 -20680 14 -20360
rect -306 -21400 14 -21080
rect -306 -22120 14 -21800
rect -306 -22840 14 -22520
<< metal4 >>
rect -198 22841 -94 23040
rect 282 22892 386 23040
rect -307 22840 15 22841
rect -307 22520 -306 22840
rect 14 22520 15 22840
rect -307 22519 15 22520
rect -198 22121 -94 22519
rect 282 22468 302 22892
rect 366 22468 386 22892
rect 282 22172 386 22468
rect -307 22120 15 22121
rect -307 21800 -306 22120
rect 14 21800 15 22120
rect -307 21799 15 21800
rect -198 21401 -94 21799
rect 282 21748 302 22172
rect 366 21748 386 22172
rect 282 21452 386 21748
rect -307 21400 15 21401
rect -307 21080 -306 21400
rect 14 21080 15 21400
rect -307 21079 15 21080
rect -198 20681 -94 21079
rect 282 21028 302 21452
rect 366 21028 386 21452
rect 282 20732 386 21028
rect -307 20680 15 20681
rect -307 20360 -306 20680
rect 14 20360 15 20680
rect -307 20359 15 20360
rect -198 19961 -94 20359
rect 282 20308 302 20732
rect 366 20308 386 20732
rect 282 20012 386 20308
rect -307 19960 15 19961
rect -307 19640 -306 19960
rect 14 19640 15 19960
rect -307 19639 15 19640
rect -198 19241 -94 19639
rect 282 19588 302 20012
rect 366 19588 386 20012
rect 282 19292 386 19588
rect -307 19240 15 19241
rect -307 18920 -306 19240
rect 14 18920 15 19240
rect -307 18919 15 18920
rect -198 18521 -94 18919
rect 282 18868 302 19292
rect 366 18868 386 19292
rect 282 18572 386 18868
rect -307 18520 15 18521
rect -307 18200 -306 18520
rect 14 18200 15 18520
rect -307 18199 15 18200
rect -198 17801 -94 18199
rect 282 18148 302 18572
rect 366 18148 386 18572
rect 282 17852 386 18148
rect -307 17800 15 17801
rect -307 17480 -306 17800
rect 14 17480 15 17800
rect -307 17479 15 17480
rect -198 17081 -94 17479
rect 282 17428 302 17852
rect 366 17428 386 17852
rect 282 17132 386 17428
rect -307 17080 15 17081
rect -307 16760 -306 17080
rect 14 16760 15 17080
rect -307 16759 15 16760
rect -198 16361 -94 16759
rect 282 16708 302 17132
rect 366 16708 386 17132
rect 282 16412 386 16708
rect -307 16360 15 16361
rect -307 16040 -306 16360
rect 14 16040 15 16360
rect -307 16039 15 16040
rect -198 15641 -94 16039
rect 282 15988 302 16412
rect 366 15988 386 16412
rect 282 15692 386 15988
rect -307 15640 15 15641
rect -307 15320 -306 15640
rect 14 15320 15 15640
rect -307 15319 15 15320
rect -198 14921 -94 15319
rect 282 15268 302 15692
rect 366 15268 386 15692
rect 282 14972 386 15268
rect -307 14920 15 14921
rect -307 14600 -306 14920
rect 14 14600 15 14920
rect -307 14599 15 14600
rect -198 14201 -94 14599
rect 282 14548 302 14972
rect 366 14548 386 14972
rect 282 14252 386 14548
rect -307 14200 15 14201
rect -307 13880 -306 14200
rect 14 13880 15 14200
rect -307 13879 15 13880
rect -198 13481 -94 13879
rect 282 13828 302 14252
rect 366 13828 386 14252
rect 282 13532 386 13828
rect -307 13480 15 13481
rect -307 13160 -306 13480
rect 14 13160 15 13480
rect -307 13159 15 13160
rect -198 12761 -94 13159
rect 282 13108 302 13532
rect 366 13108 386 13532
rect 282 12812 386 13108
rect -307 12760 15 12761
rect -307 12440 -306 12760
rect 14 12440 15 12760
rect -307 12439 15 12440
rect -198 12041 -94 12439
rect 282 12388 302 12812
rect 366 12388 386 12812
rect 282 12092 386 12388
rect -307 12040 15 12041
rect -307 11720 -306 12040
rect 14 11720 15 12040
rect -307 11719 15 11720
rect -198 11321 -94 11719
rect 282 11668 302 12092
rect 366 11668 386 12092
rect 282 11372 386 11668
rect -307 11320 15 11321
rect -307 11000 -306 11320
rect 14 11000 15 11320
rect -307 10999 15 11000
rect -198 10601 -94 10999
rect 282 10948 302 11372
rect 366 10948 386 11372
rect 282 10652 386 10948
rect -307 10600 15 10601
rect -307 10280 -306 10600
rect 14 10280 15 10600
rect -307 10279 15 10280
rect -198 9881 -94 10279
rect 282 10228 302 10652
rect 366 10228 386 10652
rect 282 9932 386 10228
rect -307 9880 15 9881
rect -307 9560 -306 9880
rect 14 9560 15 9880
rect -307 9559 15 9560
rect -198 9161 -94 9559
rect 282 9508 302 9932
rect 366 9508 386 9932
rect 282 9212 386 9508
rect -307 9160 15 9161
rect -307 8840 -306 9160
rect 14 8840 15 9160
rect -307 8839 15 8840
rect -198 8441 -94 8839
rect 282 8788 302 9212
rect 366 8788 386 9212
rect 282 8492 386 8788
rect -307 8440 15 8441
rect -307 8120 -306 8440
rect 14 8120 15 8440
rect -307 8119 15 8120
rect -198 7721 -94 8119
rect 282 8068 302 8492
rect 366 8068 386 8492
rect 282 7772 386 8068
rect -307 7720 15 7721
rect -307 7400 -306 7720
rect 14 7400 15 7720
rect -307 7399 15 7400
rect -198 7001 -94 7399
rect 282 7348 302 7772
rect 366 7348 386 7772
rect 282 7052 386 7348
rect -307 7000 15 7001
rect -307 6680 -306 7000
rect 14 6680 15 7000
rect -307 6679 15 6680
rect -198 6281 -94 6679
rect 282 6628 302 7052
rect 366 6628 386 7052
rect 282 6332 386 6628
rect -307 6280 15 6281
rect -307 5960 -306 6280
rect 14 5960 15 6280
rect -307 5959 15 5960
rect -198 5561 -94 5959
rect 282 5908 302 6332
rect 366 5908 386 6332
rect 282 5612 386 5908
rect -307 5560 15 5561
rect -307 5240 -306 5560
rect 14 5240 15 5560
rect -307 5239 15 5240
rect -198 4841 -94 5239
rect 282 5188 302 5612
rect 366 5188 386 5612
rect 282 4892 386 5188
rect -307 4840 15 4841
rect -307 4520 -306 4840
rect 14 4520 15 4840
rect -307 4519 15 4520
rect -198 4121 -94 4519
rect 282 4468 302 4892
rect 366 4468 386 4892
rect 282 4172 386 4468
rect -307 4120 15 4121
rect -307 3800 -306 4120
rect 14 3800 15 4120
rect -307 3799 15 3800
rect -198 3401 -94 3799
rect 282 3748 302 4172
rect 366 3748 386 4172
rect 282 3452 386 3748
rect -307 3400 15 3401
rect -307 3080 -306 3400
rect 14 3080 15 3400
rect -307 3079 15 3080
rect -198 2681 -94 3079
rect 282 3028 302 3452
rect 366 3028 386 3452
rect 282 2732 386 3028
rect -307 2680 15 2681
rect -307 2360 -306 2680
rect 14 2360 15 2680
rect -307 2359 15 2360
rect -198 1961 -94 2359
rect 282 2308 302 2732
rect 366 2308 386 2732
rect 282 2012 386 2308
rect -307 1960 15 1961
rect -307 1640 -306 1960
rect 14 1640 15 1960
rect -307 1639 15 1640
rect -198 1241 -94 1639
rect 282 1588 302 2012
rect 366 1588 386 2012
rect 282 1292 386 1588
rect -307 1240 15 1241
rect -307 920 -306 1240
rect 14 920 15 1240
rect -307 919 15 920
rect -198 521 -94 919
rect 282 868 302 1292
rect 366 868 386 1292
rect 282 572 386 868
rect -307 520 15 521
rect -307 200 -306 520
rect 14 200 15 520
rect -307 199 15 200
rect -198 -199 -94 199
rect 282 148 302 572
rect 366 148 386 572
rect 282 -148 386 148
rect -307 -200 15 -199
rect -307 -520 -306 -200
rect 14 -520 15 -200
rect -307 -521 15 -520
rect -198 -919 -94 -521
rect 282 -572 302 -148
rect 366 -572 386 -148
rect 282 -868 386 -572
rect -307 -920 15 -919
rect -307 -1240 -306 -920
rect 14 -1240 15 -920
rect -307 -1241 15 -1240
rect -198 -1639 -94 -1241
rect 282 -1292 302 -868
rect 366 -1292 386 -868
rect 282 -1588 386 -1292
rect -307 -1640 15 -1639
rect -307 -1960 -306 -1640
rect 14 -1960 15 -1640
rect -307 -1961 15 -1960
rect -198 -2359 -94 -1961
rect 282 -2012 302 -1588
rect 366 -2012 386 -1588
rect 282 -2308 386 -2012
rect -307 -2360 15 -2359
rect -307 -2680 -306 -2360
rect 14 -2680 15 -2360
rect -307 -2681 15 -2680
rect -198 -3079 -94 -2681
rect 282 -2732 302 -2308
rect 366 -2732 386 -2308
rect 282 -3028 386 -2732
rect -307 -3080 15 -3079
rect -307 -3400 -306 -3080
rect 14 -3400 15 -3080
rect -307 -3401 15 -3400
rect -198 -3799 -94 -3401
rect 282 -3452 302 -3028
rect 366 -3452 386 -3028
rect 282 -3748 386 -3452
rect -307 -3800 15 -3799
rect -307 -4120 -306 -3800
rect 14 -4120 15 -3800
rect -307 -4121 15 -4120
rect -198 -4519 -94 -4121
rect 282 -4172 302 -3748
rect 366 -4172 386 -3748
rect 282 -4468 386 -4172
rect -307 -4520 15 -4519
rect -307 -4840 -306 -4520
rect 14 -4840 15 -4520
rect -307 -4841 15 -4840
rect -198 -5239 -94 -4841
rect 282 -4892 302 -4468
rect 366 -4892 386 -4468
rect 282 -5188 386 -4892
rect -307 -5240 15 -5239
rect -307 -5560 -306 -5240
rect 14 -5560 15 -5240
rect -307 -5561 15 -5560
rect -198 -5959 -94 -5561
rect 282 -5612 302 -5188
rect 366 -5612 386 -5188
rect 282 -5908 386 -5612
rect -307 -5960 15 -5959
rect -307 -6280 -306 -5960
rect 14 -6280 15 -5960
rect -307 -6281 15 -6280
rect -198 -6679 -94 -6281
rect 282 -6332 302 -5908
rect 366 -6332 386 -5908
rect 282 -6628 386 -6332
rect -307 -6680 15 -6679
rect -307 -7000 -306 -6680
rect 14 -7000 15 -6680
rect -307 -7001 15 -7000
rect -198 -7399 -94 -7001
rect 282 -7052 302 -6628
rect 366 -7052 386 -6628
rect 282 -7348 386 -7052
rect -307 -7400 15 -7399
rect -307 -7720 -306 -7400
rect 14 -7720 15 -7400
rect -307 -7721 15 -7720
rect -198 -8119 -94 -7721
rect 282 -7772 302 -7348
rect 366 -7772 386 -7348
rect 282 -8068 386 -7772
rect -307 -8120 15 -8119
rect -307 -8440 -306 -8120
rect 14 -8440 15 -8120
rect -307 -8441 15 -8440
rect -198 -8839 -94 -8441
rect 282 -8492 302 -8068
rect 366 -8492 386 -8068
rect 282 -8788 386 -8492
rect -307 -8840 15 -8839
rect -307 -9160 -306 -8840
rect 14 -9160 15 -8840
rect -307 -9161 15 -9160
rect -198 -9559 -94 -9161
rect 282 -9212 302 -8788
rect 366 -9212 386 -8788
rect 282 -9508 386 -9212
rect -307 -9560 15 -9559
rect -307 -9880 -306 -9560
rect 14 -9880 15 -9560
rect -307 -9881 15 -9880
rect -198 -10279 -94 -9881
rect 282 -9932 302 -9508
rect 366 -9932 386 -9508
rect 282 -10228 386 -9932
rect -307 -10280 15 -10279
rect -307 -10600 -306 -10280
rect 14 -10600 15 -10280
rect -307 -10601 15 -10600
rect -198 -10999 -94 -10601
rect 282 -10652 302 -10228
rect 366 -10652 386 -10228
rect 282 -10948 386 -10652
rect -307 -11000 15 -10999
rect -307 -11320 -306 -11000
rect 14 -11320 15 -11000
rect -307 -11321 15 -11320
rect -198 -11719 -94 -11321
rect 282 -11372 302 -10948
rect 366 -11372 386 -10948
rect 282 -11668 386 -11372
rect -307 -11720 15 -11719
rect -307 -12040 -306 -11720
rect 14 -12040 15 -11720
rect -307 -12041 15 -12040
rect -198 -12439 -94 -12041
rect 282 -12092 302 -11668
rect 366 -12092 386 -11668
rect 282 -12388 386 -12092
rect -307 -12440 15 -12439
rect -307 -12760 -306 -12440
rect 14 -12760 15 -12440
rect -307 -12761 15 -12760
rect -198 -13159 -94 -12761
rect 282 -12812 302 -12388
rect 366 -12812 386 -12388
rect 282 -13108 386 -12812
rect -307 -13160 15 -13159
rect -307 -13480 -306 -13160
rect 14 -13480 15 -13160
rect -307 -13481 15 -13480
rect -198 -13879 -94 -13481
rect 282 -13532 302 -13108
rect 366 -13532 386 -13108
rect 282 -13828 386 -13532
rect -307 -13880 15 -13879
rect -307 -14200 -306 -13880
rect 14 -14200 15 -13880
rect -307 -14201 15 -14200
rect -198 -14599 -94 -14201
rect 282 -14252 302 -13828
rect 366 -14252 386 -13828
rect 282 -14548 386 -14252
rect -307 -14600 15 -14599
rect -307 -14920 -306 -14600
rect 14 -14920 15 -14600
rect -307 -14921 15 -14920
rect -198 -15319 -94 -14921
rect 282 -14972 302 -14548
rect 366 -14972 386 -14548
rect 282 -15268 386 -14972
rect -307 -15320 15 -15319
rect -307 -15640 -306 -15320
rect 14 -15640 15 -15320
rect -307 -15641 15 -15640
rect -198 -16039 -94 -15641
rect 282 -15692 302 -15268
rect 366 -15692 386 -15268
rect 282 -15988 386 -15692
rect -307 -16040 15 -16039
rect -307 -16360 -306 -16040
rect 14 -16360 15 -16040
rect -307 -16361 15 -16360
rect -198 -16759 -94 -16361
rect 282 -16412 302 -15988
rect 366 -16412 386 -15988
rect 282 -16708 386 -16412
rect -307 -16760 15 -16759
rect -307 -17080 -306 -16760
rect 14 -17080 15 -16760
rect -307 -17081 15 -17080
rect -198 -17479 -94 -17081
rect 282 -17132 302 -16708
rect 366 -17132 386 -16708
rect 282 -17428 386 -17132
rect -307 -17480 15 -17479
rect -307 -17800 -306 -17480
rect 14 -17800 15 -17480
rect -307 -17801 15 -17800
rect -198 -18199 -94 -17801
rect 282 -17852 302 -17428
rect 366 -17852 386 -17428
rect 282 -18148 386 -17852
rect -307 -18200 15 -18199
rect -307 -18520 -306 -18200
rect 14 -18520 15 -18200
rect -307 -18521 15 -18520
rect -198 -18919 -94 -18521
rect 282 -18572 302 -18148
rect 366 -18572 386 -18148
rect 282 -18868 386 -18572
rect -307 -18920 15 -18919
rect -307 -19240 -306 -18920
rect 14 -19240 15 -18920
rect -307 -19241 15 -19240
rect -198 -19639 -94 -19241
rect 282 -19292 302 -18868
rect 366 -19292 386 -18868
rect 282 -19588 386 -19292
rect -307 -19640 15 -19639
rect -307 -19960 -306 -19640
rect 14 -19960 15 -19640
rect -307 -19961 15 -19960
rect -198 -20359 -94 -19961
rect 282 -20012 302 -19588
rect 366 -20012 386 -19588
rect 282 -20308 386 -20012
rect -307 -20360 15 -20359
rect -307 -20680 -306 -20360
rect 14 -20680 15 -20360
rect -307 -20681 15 -20680
rect -198 -21079 -94 -20681
rect 282 -20732 302 -20308
rect 366 -20732 386 -20308
rect 282 -21028 386 -20732
rect -307 -21080 15 -21079
rect -307 -21400 -306 -21080
rect 14 -21400 15 -21080
rect -307 -21401 15 -21400
rect -198 -21799 -94 -21401
rect 282 -21452 302 -21028
rect 366 -21452 386 -21028
rect 282 -21748 386 -21452
rect -307 -21800 15 -21799
rect -307 -22120 -306 -21800
rect 14 -22120 15 -21800
rect -307 -22121 15 -22120
rect -198 -22519 -94 -22121
rect 282 -22172 302 -21748
rect 366 -22172 386 -21748
rect 282 -22468 386 -22172
rect -307 -22520 15 -22519
rect -307 -22840 -306 -22520
rect 14 -22840 15 -22520
rect -307 -22841 15 -22840
rect -198 -23040 -94 -22841
rect 282 -22892 302 -22468
rect 366 -22892 386 -22468
rect 282 -23040 386 -22892
<< properties >>
string FIXED_BBOX -386 22440 94 22920
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.0 l 2.0 val 9.52 carea 2.00 cperi 0.19 nx 1 ny 64 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
