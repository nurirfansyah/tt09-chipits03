MACRO tt_um_mbkmicdec_ringosc
  CLASS BLOCK ;
  FOREIGN tt_um_mbkmicdec_ringosc ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.000000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 120.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 120.000000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 78.010 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 78.010 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 121.335 87.745 124.435 87.845 ;
        RECT 132.665 87.745 135.765 87.845 ;
        RECT 121.335 84.425 135.765 87.745 ;
        RECT 121.335 84.155 124.435 84.425 ;
      LAYER nwell ;
        RECT 126.525 84.155 130.575 84.220 ;
      LAYER pwell ;
        RECT 132.665 84.155 135.765 84.425 ;
      LAYER nwell ;
        RECT 121.335 78.885 135.765 84.155 ;
      LAYER pwell ;
        RECT 125.780 77.610 125.950 77.635 ;
        RECT 125.780 77.465 126.880 77.610 ;
        RECT 125.970 73.740 126.880 77.465 ;
      LAYER nwell ;
        RECT 127.170 73.250 130.000 78.885 ;
      LAYER pwell ;
        RECT 131.220 77.610 131.390 77.635 ;
        RECT 130.290 77.465 131.390 77.610 ;
        RECT 130.290 73.740 131.200 77.465 ;
        RECT 114.240 23.425 118.340 73.245 ;
      LAYER nwell ;
        RECT 120.160 23.430 137.035 73.250 ;
      LAYER pwell ;
        RECT 138.855 23.425 142.955 73.245 ;
      LAYER li1 ;
        RECT 121.515 87.495 124.255 87.665 ;
        RECT 121.515 86.085 121.685 87.495 ;
        RECT 122.025 86.625 122.195 86.955 ;
        RECT 122.365 86.925 123.405 87.095 ;
        RECT 122.365 86.485 123.405 86.655 ;
        RECT 123.575 86.625 123.745 86.955 ;
        RECT 124.085 86.085 124.255 87.495 ;
        RECT 121.515 85.915 124.255 86.085 ;
        RECT 121.515 84.505 121.685 85.915 ;
        RECT 122.025 85.045 122.195 85.375 ;
        RECT 122.365 85.345 123.405 85.515 ;
        RECT 122.365 84.905 123.405 85.075 ;
        RECT 123.575 85.045 123.745 85.375 ;
        RECT 124.085 84.505 124.255 85.915 ;
        RECT 132.845 87.495 135.585 87.665 ;
        RECT 132.845 86.085 133.015 87.495 ;
        RECT 133.355 86.625 133.525 86.955 ;
        RECT 133.695 86.925 134.735 87.095 ;
        RECT 133.695 86.485 134.735 86.655 ;
        RECT 134.905 86.625 135.075 86.955 ;
        RECT 135.415 86.085 135.585 87.495 ;
        RECT 132.845 85.915 135.585 86.085 ;
        RECT 126.715 85.440 128.095 85.610 ;
        RECT 129.005 85.440 130.385 85.610 ;
        RECT 126.800 84.640 127.110 85.440 ;
        RECT 127.315 84.640 128.010 85.270 ;
        RECT 129.090 84.640 129.400 85.440 ;
        RECT 129.605 84.640 130.300 85.270 ;
        RECT 121.515 84.335 124.255 84.505 ;
        RECT 126.810 84.200 127.145 84.470 ;
        RECT 127.315 84.040 127.485 84.640 ;
        RECT 127.655 84.200 127.990 84.450 ;
        RECT 129.100 84.200 129.435 84.470 ;
        RECT 129.605 84.040 129.775 84.640 ;
        RECT 132.845 84.505 133.015 85.915 ;
        RECT 133.355 85.045 133.525 85.375 ;
        RECT 133.695 85.345 134.735 85.515 ;
        RECT 133.695 84.905 134.735 85.075 ;
        RECT 134.905 85.045 135.075 85.375 ;
        RECT 135.415 84.505 135.585 85.915 ;
        RECT 129.945 84.200 130.280 84.450 ;
        RECT 132.845 84.335 135.585 84.505 ;
        RECT 121.515 83.805 126.345 83.975 ;
        RECT 121.515 82.395 121.685 83.805 ;
        RECT 122.025 82.935 122.195 83.265 ;
        RECT 122.410 83.235 125.450 83.405 ;
        RECT 122.410 82.795 125.450 82.965 ;
        RECT 125.665 82.935 125.835 83.265 ;
        RECT 126.175 82.395 126.345 83.805 ;
        RECT 126.800 82.890 127.080 84.030 ;
        RECT 127.250 83.060 127.580 84.040 ;
        RECT 127.750 82.890 128.010 84.030 ;
        RECT 129.090 82.890 129.370 84.030 ;
        RECT 129.540 83.060 129.870 84.040 ;
        RECT 130.040 82.890 130.300 84.030 ;
        RECT 130.755 83.805 135.585 83.975 ;
        RECT 126.715 82.720 128.095 82.890 ;
        RECT 129.005 82.720 130.385 82.890 ;
        RECT 121.515 82.225 126.345 82.395 ;
        RECT 121.515 80.815 121.685 82.225 ;
        RECT 122.025 81.355 122.195 81.685 ;
        RECT 122.410 81.655 125.450 81.825 ;
        RECT 122.410 81.215 125.450 81.385 ;
        RECT 125.665 81.355 125.835 81.685 ;
        RECT 126.175 80.815 126.345 82.225 ;
        RECT 121.515 80.645 126.345 80.815 ;
        RECT 121.515 79.235 121.685 80.645 ;
        RECT 122.025 79.775 122.195 80.105 ;
        RECT 122.410 80.075 125.450 80.245 ;
        RECT 122.410 79.635 125.450 79.805 ;
        RECT 125.665 79.775 125.835 80.105 ;
        RECT 126.175 79.235 126.345 80.645 ;
        RECT 121.515 79.065 126.345 79.235 ;
        RECT 130.755 82.395 130.925 83.805 ;
        RECT 131.265 82.935 131.435 83.265 ;
        RECT 131.650 83.235 134.690 83.405 ;
        RECT 131.650 82.795 134.690 82.965 ;
        RECT 134.905 82.935 135.075 83.265 ;
        RECT 135.415 82.395 135.585 83.805 ;
        RECT 130.755 82.225 135.585 82.395 ;
        RECT 130.755 80.815 130.925 82.225 ;
        RECT 131.265 81.355 131.435 81.685 ;
        RECT 131.650 81.655 134.690 81.825 ;
        RECT 131.650 81.215 134.690 81.385 ;
        RECT 134.905 81.355 135.075 81.685 ;
        RECT 135.415 80.815 135.585 82.225 ;
        RECT 130.755 80.645 135.585 80.815 ;
        RECT 130.755 79.235 130.925 80.645 ;
        RECT 131.265 79.775 131.435 80.105 ;
        RECT 131.650 80.075 134.690 80.245 ;
        RECT 131.650 79.635 134.690 79.805 ;
        RECT 134.905 79.775 135.075 80.105 ;
        RECT 135.415 79.235 135.585 80.645 ;
        RECT 130.755 79.065 135.585 79.235 ;
        RECT 125.780 77.525 125.950 77.780 ;
        RECT 125.780 77.270 126.410 77.525 ;
        RECT 126.580 77.350 127.530 77.695 ;
        RECT 128.500 77.525 128.670 77.780 ;
        RECT 125.780 76.600 125.950 77.270 ;
        RECT 126.580 77.100 126.770 77.350 ;
        RECT 127.360 77.100 127.530 77.350 ;
        RECT 127.700 77.270 129.470 77.525 ;
        RECT 129.640 77.350 130.590 77.695 ;
        RECT 131.220 77.525 131.390 77.780 ;
        RECT 126.120 76.770 126.770 77.100 ;
        RECT 125.780 76.430 126.410 76.600 ;
        RECT 125.780 75.760 125.950 76.430 ;
        RECT 126.580 76.260 126.770 76.770 ;
        RECT 126.120 75.930 126.770 76.260 ;
        RECT 125.780 75.590 126.410 75.760 ;
        RECT 125.780 74.920 125.950 75.590 ;
        RECT 126.580 75.420 126.770 75.930 ;
        RECT 126.120 75.090 126.770 75.420 ;
        RECT 125.780 74.750 126.410 74.920 ;
        RECT 125.780 74.080 125.950 74.750 ;
        RECT 126.580 74.580 126.770 75.090 ;
        RECT 126.120 74.250 126.770 74.580 ;
        RECT 125.780 73.775 126.410 74.080 ;
        RECT 126.580 74.045 126.770 74.250 ;
        RECT 126.940 74.245 127.190 77.100 ;
        RECT 127.360 76.770 128.330 77.100 ;
        RECT 127.360 76.260 127.530 76.770 ;
        RECT 128.500 76.600 128.670 77.270 ;
        RECT 129.640 77.100 129.810 77.350 ;
        RECT 130.400 77.100 130.590 77.350 ;
        RECT 130.760 77.270 131.390 77.525 ;
        RECT 128.840 76.770 129.810 77.100 ;
        RECT 127.700 76.430 129.470 76.600 ;
        RECT 127.360 75.930 128.330 76.260 ;
        RECT 127.360 75.420 127.530 75.930 ;
        RECT 128.500 75.760 128.670 76.430 ;
        RECT 129.640 76.260 129.810 76.770 ;
        RECT 128.840 75.930 129.810 76.260 ;
        RECT 127.700 75.590 129.470 75.760 ;
        RECT 127.360 75.090 128.330 75.420 ;
        RECT 127.360 74.580 127.530 75.090 ;
        RECT 128.500 74.920 128.670 75.590 ;
        RECT 129.640 75.420 129.810 75.930 ;
        RECT 128.840 75.090 129.810 75.420 ;
        RECT 127.700 74.750 129.470 74.920 ;
        RECT 127.360 74.250 128.330 74.580 ;
        RECT 126.940 74.215 127.110 74.245 ;
        RECT 127.360 74.045 127.530 74.250 ;
        RECT 128.500 74.080 128.670 74.750 ;
        RECT 129.640 74.580 129.810 75.090 ;
        RECT 128.840 74.250 129.810 74.580 ;
        RECT 125.780 73.640 125.950 73.775 ;
        RECT 126.580 73.725 127.530 74.045 ;
        RECT 127.700 73.780 129.470 74.080 ;
        RECT 129.640 74.045 129.810 74.250 ;
        RECT 129.980 74.245 130.230 77.100 ;
        RECT 130.400 76.770 131.050 77.100 ;
        RECT 130.400 76.260 130.590 76.770 ;
        RECT 131.220 76.600 131.390 77.270 ;
        RECT 130.760 76.430 131.390 76.600 ;
        RECT 130.400 75.930 131.050 76.260 ;
        RECT 130.400 75.420 130.590 75.930 ;
        RECT 131.220 75.760 131.390 76.430 ;
        RECT 130.760 75.590 131.390 75.760 ;
        RECT 130.400 75.090 131.050 75.420 ;
        RECT 130.400 74.580 130.590 75.090 ;
        RECT 131.220 74.920 131.390 75.590 ;
        RECT 130.760 74.750 131.390 74.920 ;
        RECT 130.400 74.250 131.050 74.580 ;
        RECT 130.400 74.045 130.590 74.250 ;
        RECT 131.220 74.080 131.390 74.750 ;
        RECT 128.500 73.640 128.670 73.780 ;
        RECT 129.640 73.725 130.590 74.045 ;
        RECT 130.760 73.775 131.390 74.080 ;
        RECT 131.220 73.640 131.390 73.775 ;
        RECT 113.740 73.245 114.240 73.425 ;
        RECT 113.740 72.895 118.160 73.245 ;
        RECT 113.740 56.635 114.590 72.895 ;
        RECT 115.270 72.325 117.310 72.495 ;
        RECT 114.930 57.265 115.100 72.265 ;
        RECT 117.480 57.265 117.650 72.265 ;
        RECT 115.270 57.035 117.310 57.205 ;
        RECT 117.990 56.635 118.160 72.895 ;
        RECT 113.740 56.465 118.160 56.635 ;
        RECT 113.740 40.205 114.590 56.465 ;
        RECT 115.270 55.895 117.310 56.065 ;
        RECT 114.930 40.835 115.100 55.835 ;
        RECT 117.480 40.835 117.650 55.835 ;
        RECT 115.270 40.605 117.310 40.775 ;
        RECT 117.990 40.205 118.160 56.465 ;
        RECT 113.740 40.035 118.160 40.205 ;
        RECT 113.740 23.775 114.590 40.035 ;
        RECT 115.270 39.465 117.310 39.635 ;
        RECT 114.930 24.405 115.100 39.405 ;
        RECT 117.480 24.405 117.650 39.405 ;
        RECT 115.270 24.175 117.310 24.345 ;
        RECT 117.990 23.775 118.160 40.035 ;
        RECT 113.740 23.425 118.160 23.775 ;
        RECT 120.340 72.900 128.350 73.250 ;
        RECT 120.340 56.640 120.510 72.900 ;
        RECT 121.235 72.330 127.275 72.500 ;
        RECT 120.850 57.270 121.020 72.270 ;
        RECT 127.490 57.270 127.660 72.270 ;
        RECT 121.235 57.040 127.275 57.210 ;
        RECT 128.000 56.640 128.350 72.900 ;
        RECT 120.340 56.470 128.350 56.640 ;
        RECT 120.340 40.210 120.510 56.470 ;
        RECT 121.235 55.900 127.275 56.070 ;
        RECT 120.850 40.840 121.020 55.840 ;
        RECT 127.490 40.840 127.660 55.840 ;
        RECT 121.235 40.610 127.275 40.780 ;
        RECT 128.000 40.210 128.350 56.470 ;
        RECT 120.340 40.040 128.350 40.210 ;
        RECT 120.340 23.780 120.510 40.040 ;
        RECT 121.235 39.470 127.275 39.640 ;
        RECT 120.850 24.410 121.020 39.410 ;
        RECT 127.490 24.410 127.660 39.410 ;
        RECT 121.235 24.180 127.275 24.350 ;
        RECT 128.000 23.780 128.350 40.040 ;
        RECT 120.340 23.430 128.350 23.780 ;
        RECT 128.845 72.900 136.855 73.250 ;
        RECT 142.955 73.245 143.455 73.425 ;
        RECT 128.845 56.640 129.195 72.900 ;
        RECT 129.920 72.330 135.960 72.500 ;
        RECT 129.535 57.270 129.705 72.270 ;
        RECT 136.175 57.270 136.345 72.270 ;
        RECT 129.920 57.040 135.960 57.210 ;
        RECT 136.685 56.640 136.855 72.900 ;
        RECT 128.845 56.470 136.855 56.640 ;
        RECT 128.845 40.210 129.195 56.470 ;
        RECT 129.920 55.900 135.960 56.070 ;
        RECT 129.535 40.840 129.705 55.840 ;
        RECT 136.175 40.840 136.345 55.840 ;
        RECT 129.920 40.610 135.960 40.780 ;
        RECT 136.685 40.210 136.855 56.470 ;
        RECT 128.845 40.040 136.855 40.210 ;
        RECT 128.845 23.780 129.195 40.040 ;
        RECT 129.920 39.470 135.960 39.640 ;
        RECT 129.535 24.410 129.705 39.410 ;
        RECT 136.175 24.410 136.345 39.410 ;
        RECT 129.920 24.180 135.960 24.350 ;
        RECT 136.685 23.780 136.855 40.040 ;
        RECT 128.845 23.430 136.855 23.780 ;
        RECT 139.035 72.895 143.455 73.245 ;
        RECT 139.035 56.635 139.205 72.895 ;
        RECT 139.885 72.325 141.925 72.495 ;
        RECT 139.545 57.265 139.715 72.265 ;
        RECT 142.095 57.265 142.265 72.265 ;
        RECT 139.885 57.035 141.925 57.205 ;
        RECT 142.605 56.635 143.455 72.895 ;
        RECT 139.035 56.465 143.455 56.635 ;
        RECT 139.035 40.205 139.205 56.465 ;
        RECT 139.885 55.895 141.925 56.065 ;
        RECT 139.545 40.835 139.715 55.835 ;
        RECT 142.095 40.835 142.265 55.835 ;
        RECT 139.885 40.605 141.925 40.775 ;
        RECT 142.605 40.205 143.455 56.465 ;
        RECT 139.035 40.035 143.455 40.205 ;
        RECT 139.035 23.775 139.205 40.035 ;
        RECT 139.885 39.465 141.925 39.635 ;
        RECT 139.545 24.405 139.715 39.405 ;
        RECT 142.095 24.405 142.265 39.405 ;
        RECT 139.885 24.175 141.925 24.345 ;
        RECT 142.605 23.775 143.455 40.035 ;
        RECT 139.035 23.425 143.455 23.775 ;
      LAYER met1 ;
        RECT 113.190 87.845 115.290 88.570 ;
        RECT 113.190 87.360 143.485 87.845 ;
        RECT 113.190 86.570 115.290 87.360 ;
        RECT 123.135 87.125 123.385 87.360 ;
        RECT 121.285 86.625 121.665 86.955 ;
        RECT 121.845 86.625 122.225 86.955 ;
        RECT 122.385 86.895 123.385 87.125 ;
        RECT 113.710 77.560 114.270 86.570 ;
        RECT 121.335 81.685 121.595 86.625 ;
        RECT 122.385 86.455 123.385 86.685 ;
        RECT 123.545 86.625 123.825 86.955 ;
        RECT 123.135 85.545 123.385 86.455 ;
        RECT 130.070 85.765 130.385 87.360 ;
        RECT 133.715 87.125 133.965 87.360 ;
        RECT 133.275 86.625 133.555 86.955 ;
        RECT 133.715 86.895 134.715 87.125 ;
        RECT 133.715 86.455 134.715 86.685 ;
        RECT 134.875 86.625 135.255 86.955 ;
        RECT 135.435 86.625 135.815 86.955 ;
        RECT 121.945 84.595 122.225 85.375 ;
        RECT 122.385 85.315 123.385 85.545 ;
        RECT 122.385 84.875 123.385 85.105 ;
        RECT 123.545 85.045 123.825 85.375 ;
        RECT 126.715 85.285 130.390 85.765 ;
        RECT 133.715 85.545 133.965 86.455 ;
        RECT 121.895 84.335 122.275 84.595 ;
        RECT 121.945 82.935 122.225 84.335 ;
        RECT 123.135 83.975 123.385 84.875 ;
        RECT 127.640 84.810 128.675 85.090 ;
        RECT 129.720 84.835 130.110 85.115 ;
        RECT 133.275 85.045 133.555 85.375 ;
        RECT 133.715 85.315 134.715 85.545 ;
        RECT 133.715 84.875 134.715 85.105 ;
        RECT 126.800 84.135 127.135 84.480 ;
        RECT 123.085 83.715 123.465 83.975 ;
        RECT 126.165 83.715 126.525 83.975 ;
        RECT 126.750 83.865 127.185 84.135 ;
        RECT 123.135 83.435 123.385 83.715 ;
        RECT 122.430 83.205 125.430 83.435 ;
        RECT 122.430 82.765 125.480 82.995 ;
        RECT 125.635 82.935 125.915 83.265 ;
        RECT 125.120 82.735 125.480 82.765 ;
        RECT 126.215 82.395 126.475 83.715 ;
        RECT 127.655 83.695 127.990 84.530 ;
        RECT 128.395 84.505 128.675 84.810 ;
        RECT 133.715 84.595 133.965 84.875 ;
        RECT 128.395 84.225 129.435 84.505 ;
        RECT 129.895 84.200 130.330 84.530 ;
        RECT 130.575 84.335 130.935 84.595 ;
        RECT 133.635 84.335 134.015 84.595 ;
        RECT 127.655 83.525 129.850 83.695 ;
        RECT 127.655 83.360 129.900 83.525 ;
        RECT 129.510 83.245 129.900 83.360 ;
        RECT 126.715 82.565 130.385 83.045 ;
        RECT 125.120 82.135 125.480 82.395 ;
        RECT 126.165 82.135 126.525 82.395 ;
        RECT 125.170 81.855 125.430 82.135 ;
        RECT 121.285 81.355 121.665 81.685 ;
        RECT 121.895 81.355 122.275 81.685 ;
        RECT 122.430 81.625 125.430 81.855 ;
        RECT 125.170 81.620 125.430 81.625 ;
        RECT 122.430 81.185 125.430 81.415 ;
        RECT 125.585 81.355 125.965 81.685 ;
        RECT 122.430 80.275 122.680 81.185 ;
        RECT 125.585 80.465 125.965 80.795 ;
        RECT 121.895 79.775 122.275 80.105 ;
        RECT 122.430 80.045 125.430 80.275 ;
        RECT 125.635 80.105 125.915 80.465 ;
        RECT 122.430 79.605 125.430 79.835 ;
        RECT 125.585 79.775 125.965 80.105 ;
        RECT 125.180 79.370 125.430 79.605 ;
        RECT 128.295 79.370 128.895 79.405 ;
        RECT 130.070 79.370 130.385 82.565 ;
        RECT 130.625 82.395 130.885 84.335 ;
        RECT 133.715 83.435 133.965 84.335 ;
        RECT 134.875 83.975 135.155 85.375 ;
        RECT 134.825 83.715 135.205 83.975 ;
        RECT 131.185 82.935 131.465 83.265 ;
        RECT 131.670 83.205 134.670 83.435 ;
        RECT 131.620 82.765 134.670 82.995 ;
        RECT 134.875 82.935 135.155 83.715 ;
        RECT 131.620 82.735 131.980 82.765 ;
        RECT 130.575 82.135 130.935 82.395 ;
        RECT 131.620 82.135 131.980 82.395 ;
        RECT 131.670 81.855 131.930 82.135 ;
        RECT 130.525 81.355 130.905 81.685 ;
        RECT 131.135 81.355 131.515 81.685 ;
        RECT 131.670 81.625 134.670 81.855 ;
        RECT 135.505 81.685 135.765 86.625 ;
        RECT 130.575 80.795 130.855 81.355 ;
        RECT 131.670 81.185 134.670 81.415 ;
        RECT 134.825 81.355 135.205 81.685 ;
        RECT 135.435 81.355 135.815 81.685 ;
        RECT 130.575 80.465 130.975 80.795 ;
        RECT 130.575 80.415 130.855 80.465 ;
        RECT 134.420 80.275 134.670 81.185 ;
        RECT 131.135 79.775 131.515 80.105 ;
        RECT 131.670 80.045 134.670 80.275 ;
        RECT 131.670 79.605 134.670 79.835 ;
        RECT 134.875 79.775 135.155 80.105 ;
        RECT 131.670 79.370 131.920 79.605 ;
        RECT 121.335 78.885 135.765 79.370 ;
        RECT 125.625 77.560 126.105 77.780 ;
        RECT 113.710 77.060 126.105 77.560 ;
        RECT 126.890 77.300 127.200 77.745 ;
        RECT 113.710 40.545 114.270 77.060 ;
        RECT 125.625 73.640 126.105 77.060 ;
        RECT 119.660 72.765 120.160 73.065 ;
        RECT 126.910 72.765 127.140 76.860 ;
        RECT 115.290 72.515 127.255 72.765 ;
        RECT 128.295 72.650 128.895 78.885 ;
        RECT 129.945 77.300 130.255 77.745 ;
        RECT 131.065 77.555 131.545 77.780 ;
        RECT 142.925 77.555 143.485 87.360 ;
        RECT 131.065 77.055 143.485 77.555 ;
        RECT 130.030 72.765 130.260 76.860 ;
        RECT 131.065 73.640 131.545 77.055 ;
        RECT 137.035 72.765 137.535 73.065 ;
        RECT 115.290 72.265 117.290 72.515 ;
        RECT 119.660 72.465 120.160 72.515 ;
        RECT 121.255 72.270 127.255 72.515 ;
        RECT 114.900 57.285 115.130 72.245 ;
        RECT 117.450 57.535 117.680 72.245 ;
        RECT 119.575 57.535 120.235 57.610 ;
        RECT 120.820 57.535 121.050 72.250 ;
        RECT 115.290 56.925 117.290 57.315 ;
        RECT 117.450 57.285 121.050 57.535 ;
        RECT 127.460 57.290 127.690 72.250 ;
        RECT 119.575 57.010 120.235 57.285 ;
        RECT 121.255 56.980 127.255 57.240 ;
        RECT 128.140 56.980 129.055 72.650 ;
        RECT 129.940 72.515 141.905 72.765 ;
        RECT 129.940 72.270 135.940 72.515 ;
        RECT 137.035 72.465 137.535 72.515 ;
        RECT 139.905 72.265 141.905 72.515 ;
        RECT 129.505 57.290 129.735 72.250 ;
        RECT 136.145 57.535 136.375 72.250 ;
        RECT 136.960 57.535 137.620 57.610 ;
        RECT 139.515 57.535 139.745 72.245 ;
        RECT 136.145 57.285 139.745 57.535 ;
        RECT 129.940 56.980 135.940 57.240 ;
        RECT 136.960 57.010 137.620 57.285 ;
        RECT 121.255 56.670 135.940 56.980 ;
        RECT 139.905 56.925 141.905 57.315 ;
        RECT 142.065 57.285 142.295 72.245 ;
        RECT 120.760 56.440 136.435 56.670 ;
        RECT 114.630 55.815 114.930 55.885 ;
        RECT 114.630 40.855 115.130 55.815 ;
        RECT 115.290 55.785 117.290 56.175 ;
        RECT 121.255 56.130 135.940 56.440 ;
        RECT 121.255 55.870 127.255 56.130 ;
        RECT 127.660 55.820 127.960 55.890 ;
        RECT 117.450 40.855 117.680 55.815 ;
        RECT 120.820 40.860 121.050 55.820 ;
        RECT 114.630 40.785 114.930 40.855 ;
        RECT 115.290 40.545 117.290 40.805 ;
        RECT 113.710 39.695 117.290 40.545 ;
        RECT 121.255 40.500 127.255 40.890 ;
        RECT 127.460 40.860 127.960 55.820 ;
        RECT 127.660 40.790 127.960 40.860 ;
        RECT 128.140 40.460 129.055 56.130 ;
        RECT 129.235 55.820 129.535 55.890 ;
        RECT 129.940 55.870 135.940 56.130 ;
        RECT 129.235 40.860 129.735 55.820 ;
        RECT 129.235 40.790 129.535 40.860 ;
        RECT 129.940 40.500 135.940 40.890 ;
        RECT 136.145 40.860 136.375 55.820 ;
        RECT 139.515 40.855 139.745 55.815 ;
        RECT 139.905 55.785 141.905 56.175 ;
        RECT 142.265 55.815 142.565 55.885 ;
        RECT 142.065 40.855 142.565 55.815 ;
        RECT 139.905 40.545 141.905 40.805 ;
        RECT 142.265 40.785 142.565 40.855 ;
        RECT 142.925 40.545 143.485 77.055 ;
        RECT 128.295 39.790 128.895 40.460 ;
        RECT 113.710 23.365 114.270 39.695 ;
        RECT 115.290 39.435 117.290 39.695 ;
        RECT 114.900 24.425 115.130 39.385 ;
        RECT 117.450 24.675 117.680 39.385 ;
        RECT 118.340 24.675 118.840 24.975 ;
        RECT 120.820 24.675 121.050 39.390 ;
        RECT 121.255 39.360 127.255 39.750 ;
        RECT 117.450 24.425 121.050 24.675 ;
        RECT 127.460 24.430 127.690 39.390 ;
        RECT 115.290 24.155 117.290 24.405 ;
        RECT 118.340 24.375 118.840 24.425 ;
        RECT 121.255 24.155 127.255 24.410 ;
        RECT 115.290 23.905 127.255 24.155 ;
        RECT 128.140 24.030 129.055 39.790 ;
        RECT 129.505 24.430 129.735 39.390 ;
        RECT 129.940 39.360 135.940 39.750 ;
        RECT 139.905 39.695 143.485 40.545 ;
        RECT 139.905 39.435 141.905 39.695 ;
        RECT 136.145 24.675 136.375 39.390 ;
        RECT 138.355 24.675 138.855 24.975 ;
        RECT 139.515 24.675 139.745 39.385 ;
        RECT 136.145 24.425 139.745 24.675 ;
        RECT 142.065 24.425 142.295 39.385 ;
        RECT 129.940 24.155 135.940 24.410 ;
        RECT 138.355 24.375 138.855 24.425 ;
        RECT 139.905 24.155 141.905 24.405 ;
        RECT 119.660 23.605 120.160 23.905 ;
        RECT 128.295 23.370 128.895 24.030 ;
        RECT 129.940 23.905 141.905 24.155 ;
        RECT 137.035 23.605 137.535 23.905 ;
        RECT 142.925 23.365 143.485 39.695 ;
        RECT 127.610 22.925 128.010 22.975 ;
        RECT 142.215 22.925 142.615 22.975 ;
        RECT 127.610 22.525 142.615 22.925 ;
        RECT 127.610 22.475 128.010 22.525 ;
        RECT 142.215 22.475 142.615 22.525 ;
        RECT 114.580 21.945 114.980 21.995 ;
        RECT 129.185 21.945 129.585 21.995 ;
        RECT 114.580 21.545 129.585 21.945 ;
        RECT 114.580 21.495 114.980 21.545 ;
        RECT 129.185 21.495 129.585 21.545 ;
        RECT 118.290 20.730 118.890 20.780 ;
        RECT 129.930 20.730 130.330 20.780 ;
        RECT 138.305 20.730 138.905 20.780 ;
        RECT 118.290 20.130 138.905 20.730 ;
        RECT 118.290 20.080 118.890 20.130 ;
        RECT 129.930 20.080 130.330 20.130 ;
        RECT 138.305 20.080 138.905 20.130 ;
      LAYER met2 ;
        RECT 125.760 88.995 126.020 89.255 ;
        RECT 131.145 89.245 131.425 89.255 ;
        RECT 113.240 86.520 115.240 88.620 ;
        RECT 125.675 88.410 126.170 88.995 ;
        RECT 131.045 88.660 131.540 89.245 ;
        RECT 121.335 86.955 121.615 87.005 ;
        RECT 121.895 86.955 122.175 87.005 ;
        RECT 121.335 86.625 122.175 86.955 ;
        RECT 121.335 86.575 121.615 86.625 ;
        RECT 121.895 86.575 122.175 86.625 ;
        RECT 125.760 85.070 126.020 88.410 ;
        RECT 127.690 85.070 127.980 85.140 ;
        RECT 125.760 84.810 127.980 85.070 ;
        RECT 127.690 84.760 127.980 84.810 ;
        RECT 129.770 85.115 130.060 85.165 ;
        RECT 131.145 85.115 131.425 88.660 ;
        RECT 134.925 86.955 135.205 87.005 ;
        RECT 135.485 86.955 135.765 87.005 ;
        RECT 134.925 86.625 135.765 86.955 ;
        RECT 134.925 86.575 135.205 86.625 ;
        RECT 135.485 86.575 135.765 86.625 ;
        RECT 129.770 84.835 131.425 85.115 ;
        RECT 129.770 84.785 130.060 84.835 ;
        RECT 121.945 84.595 122.225 84.645 ;
        RECT 130.625 84.595 130.885 84.645 ;
        RECT 133.685 84.595 133.965 84.645 ;
        RECT 121.945 84.335 133.965 84.595 ;
        RECT 121.945 84.285 122.225 84.335 ;
        RECT 123.135 83.975 123.415 84.025 ;
        RECT 126.215 83.975 126.475 84.025 ;
        RECT 126.800 83.975 127.135 84.185 ;
        RECT 129.945 84.150 130.280 84.335 ;
        RECT 130.625 84.285 130.885 84.335 ;
        RECT 133.685 84.285 133.965 84.335 ;
        RECT 134.875 83.975 135.155 84.025 ;
        RECT 123.135 83.715 135.155 83.975 ;
        RECT 123.135 83.665 123.415 83.715 ;
        RECT 126.215 83.665 126.475 83.715 ;
        RECT 134.875 83.665 135.155 83.715 ;
        RECT 129.560 83.195 129.850 83.575 ;
        RECT 125.170 82.995 125.430 83.045 ;
        RECT 131.670 82.995 131.930 83.045 ;
        RECT 125.170 82.735 131.930 82.995 ;
        RECT 125.170 82.685 125.430 82.735 ;
        RECT 126.845 82.515 127.105 82.735 ;
        RECT 127.770 82.515 128.030 82.735 ;
        RECT 129.150 82.515 129.410 82.735 ;
        RECT 130.070 82.515 130.330 82.735 ;
        RECT 131.670 82.685 131.930 82.735 ;
        RECT 125.170 82.395 125.430 82.445 ;
        RECT 126.215 82.395 126.475 82.445 ;
        RECT 125.170 82.135 126.475 82.395 ;
        RECT 125.170 82.085 125.430 82.135 ;
        RECT 126.215 82.085 126.475 82.135 ;
        RECT 130.625 82.395 130.885 82.445 ;
        RECT 131.670 82.395 131.930 82.445 ;
        RECT 130.625 82.135 131.930 82.395 ;
        RECT 130.625 82.085 130.885 82.135 ;
        RECT 131.670 82.085 131.930 82.135 ;
        RECT 121.335 81.685 121.615 81.735 ;
        RECT 121.945 81.685 122.225 81.735 ;
        RECT 121.335 81.355 122.225 81.685 ;
        RECT 121.335 81.305 121.615 81.355 ;
        RECT 121.945 81.305 122.225 81.355 ;
        RECT 125.635 81.685 125.915 81.735 ;
        RECT 126.245 81.685 126.525 81.735 ;
        RECT 125.635 81.355 126.525 81.685 ;
        RECT 125.635 81.305 125.915 81.355 ;
        RECT 126.245 81.305 126.525 81.355 ;
        RECT 130.575 81.685 130.855 81.735 ;
        RECT 131.185 81.685 131.465 81.735 ;
        RECT 130.575 81.355 131.465 81.685 ;
        RECT 130.575 81.305 130.855 81.355 ;
        RECT 131.185 81.305 131.465 81.355 ;
        RECT 134.875 81.685 135.155 81.735 ;
        RECT 135.485 81.685 135.765 81.735 ;
        RECT 134.875 81.355 135.765 81.685 ;
        RECT 134.875 81.305 135.155 81.355 ;
        RECT 135.485 81.305 135.765 81.355 ;
        RECT 1.000 81.130 3.000 81.180 ;
        RECT 1.000 79.130 111.930 81.130 ;
        RECT 125.635 80.795 125.915 80.845 ;
        RECT 130.640 80.795 130.925 80.845 ;
        RECT 125.635 80.465 130.925 80.795 ;
        RECT 125.635 80.415 125.915 80.465 ;
        RECT 121.945 80.105 122.225 80.155 ;
        RECT 121.335 79.775 122.225 80.105 ;
        RECT 121.945 79.725 122.225 79.775 ;
        RECT 125.635 79.725 125.915 80.155 ;
        RECT 126.915 80.080 127.170 80.160 ;
        RECT 126.855 79.800 127.235 80.080 ;
        RECT 1.000 79.080 3.000 79.130 ;
        RECT 110.450 11.500 110.925 79.130 ;
        RECT 126.915 77.695 127.170 79.800 ;
        RECT 126.840 77.350 127.250 77.695 ;
        RECT 119.610 72.515 120.210 73.250 ;
        RECT 119.605 57.535 120.205 57.640 ;
        RECT 115.240 55.835 117.340 57.265 ;
        RECT 119.605 57.040 120.210 57.535 ;
        RECT 114.580 21.945 114.980 55.835 ;
        RECT 114.530 21.545 115.030 21.945 ;
        RECT 118.290 20.730 118.890 24.925 ;
        RECT 119.605 24.155 120.205 57.040 ;
        RECT 121.205 39.410 127.305 40.840 ;
        RECT 119.605 23.655 120.210 24.155 ;
        RECT 119.605 23.650 120.205 23.655 ;
        RECT 127.610 22.925 128.010 55.840 ;
        RECT 127.560 22.525 128.060 22.925 ;
        RECT 128.320 22.765 128.880 79.400 ;
        RECT 129.970 77.695 130.230 80.465 ;
        RECT 130.640 80.415 130.925 80.465 ;
        RECT 131.185 79.725 131.465 80.155 ;
        RECT 129.895 77.350 130.305 77.695 ;
        RECT 136.985 72.515 137.585 73.250 ;
        RECT 136.990 57.535 137.590 57.640 ;
        RECT 136.985 57.040 137.590 57.535 ;
        RECT 118.240 20.130 118.940 20.730 ;
        RECT 127.610 19.025 128.010 22.525 ;
        RECT 127.550 18.470 128.060 19.025 ;
        RECT 128.360 11.500 128.835 22.765 ;
        RECT 129.185 21.945 129.585 55.840 ;
        RECT 129.890 39.410 135.990 40.840 ;
        RECT 136.990 24.155 137.590 57.040 ;
        RECT 139.855 55.835 141.955 57.265 ;
        RECT 136.985 23.655 137.590 24.155 ;
        RECT 136.990 23.650 137.590 23.655 ;
        RECT 129.135 21.545 129.635 21.945 ;
        RECT 129.185 19.025 129.585 21.545 ;
        RECT 138.305 20.780 138.905 24.925 ;
        RECT 142.215 22.925 142.615 55.835 ;
        RECT 142.165 22.525 142.665 22.925 ;
        RECT 138.300 20.730 138.910 20.780 ;
        RECT 129.880 20.130 130.380 20.730 ;
        RECT 138.255 20.130 138.955 20.730 ;
        RECT 129.130 18.470 129.640 19.025 ;
        RECT 129.930 18.520 130.330 20.130 ;
        RECT 138.300 20.080 138.910 20.130 ;
        RECT 110.450 11.025 128.835 11.500 ;
      LAYER met3 ;
        RECT 113.190 86.545 115.290 88.595 ;
        RECT 125.625 88.435 126.220 88.970 ;
        RECT 130.995 88.685 131.590 89.220 ;
        RECT 0.950 79.105 3.050 81.155 ;
        RECT 126.195 80.155 126.575 81.710 ;
        RECT 126.145 80.130 126.625 80.155 ;
        RECT 126.145 79.750 127.210 80.130 ;
        RECT 126.145 79.725 126.625 79.750 ;
        RECT 131.085 79.670 131.565 80.205 ;
        RECT 138.250 20.105 138.960 20.755 ;
        RECT 127.500 18.495 128.110 19.000 ;
        RECT 129.080 18.495 129.690 19.000 ;
      LAYER met4 ;
        RECT 1.000 81.135 3.000 220.760 ;
        RECT 4.000 88.570 6.000 220.760 ;
        RECT 91.390 91.865 91.690 224.760 ;
        RECT 94.150 94.065 94.450 224.760 ;
        RECT 94.150 93.765 131.445 94.065 ;
        RECT 91.390 91.565 126.070 91.865 ;
        RECT 125.770 88.950 126.070 91.565 ;
        RECT 131.145 89.200 131.445 93.765 ;
        RECT 113.235 88.570 115.245 88.575 ;
        RECT 4.000 86.570 115.245 88.570 ;
        RECT 125.670 88.455 126.175 88.950 ;
        RECT 131.040 88.705 131.545 89.200 ;
        RECT 0.995 79.125 3.005 81.135 ;
        RECT 1.000 78.010 3.000 79.125 ;
        RECT 4.000 78.010 6.000 86.570 ;
        RECT 113.235 86.565 115.245 86.570 ;
        RECT 126.190 79.720 131.520 80.160 ;
        RECT 138.295 20.525 138.915 20.735 ;
        RECT 143.830 20.525 144.130 224.760 ;
        RECT 138.295 20.225 144.130 20.525 ;
        RECT 138.295 20.125 138.915 20.225 ;
        RECT 127.350 13.530 128.250 19.270 ;
        RECT 128.945 15.410 129.845 19.255 ;
        RECT 128.945 14.510 152.710 15.410 ;
        RECT 127.350 12.630 133.390 13.530 ;
        RECT 132.490 1.000 133.390 12.630 ;
        RECT 151.810 1.000 152.710 14.510 ;
  END
END tt_um_mbkmicdec_ringosc
END LIBRARY

