magic
tech sky130A
magscale 1 2
timestamp 1730568870
<< error_p >>
rect -29 599 29 605
rect -29 565 -17 599
rect -29 559 29 565
rect -29 389 29 395
rect -29 355 -17 389
rect -29 349 29 355
rect -29 281 29 287
rect -29 247 -17 281
rect -29 241 29 247
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -247 29 -241
rect -29 -281 -17 -247
rect -29 -287 29 -281
rect -29 -355 29 -349
rect -29 -389 -17 -355
rect -29 -395 29 -389
rect -29 -565 29 -559
rect -29 -599 -17 -565
rect -29 -605 29 -599
<< pwell >>
rect -226 -737 226 737
<< nmos >>
rect -30 427 30 527
rect -30 109 30 209
rect -30 -209 30 -109
rect -30 -527 30 -427
<< ndiff >>
rect -88 515 -30 527
rect -88 439 -76 515
rect -42 439 -30 515
rect -88 427 -30 439
rect 30 515 88 527
rect 30 439 42 515
rect 76 439 88 515
rect 30 427 88 439
rect -88 197 -30 209
rect -88 121 -76 197
rect -42 121 -30 197
rect -88 109 -30 121
rect 30 197 88 209
rect 30 121 42 197
rect 76 121 88 197
rect 30 109 88 121
rect -88 -121 -30 -109
rect -88 -197 -76 -121
rect -42 -197 -30 -121
rect -88 -209 -30 -197
rect 30 -121 88 -109
rect 30 -197 42 -121
rect 76 -197 88 -121
rect 30 -209 88 -197
rect -88 -439 -30 -427
rect -88 -515 -76 -439
rect -42 -515 -30 -439
rect -88 -527 -30 -515
rect 30 -439 88 -427
rect 30 -515 42 -439
rect 76 -515 88 -439
rect 30 -527 88 -515
<< ndiffc >>
rect -76 439 -42 515
rect 42 439 76 515
rect -76 121 -42 197
rect 42 121 76 197
rect -76 -197 -42 -121
rect 42 -197 76 -121
rect -76 -515 -42 -439
rect 42 -515 76 -439
<< psubdiff >>
rect -190 667 -94 701
rect 94 667 190 701
rect -190 605 -156 667
rect 156 605 190 667
rect -190 -667 -156 -605
rect 156 -667 190 -605
rect -190 -701 -94 -667
rect 94 -701 190 -667
<< psubdiffcont >>
rect -94 667 94 701
rect -190 -605 -156 605
rect 156 -605 190 605
rect -94 -701 94 -667
<< poly >>
rect -33 599 33 615
rect -33 565 -17 599
rect 17 565 33 599
rect -33 549 33 565
rect -30 527 30 549
rect -30 405 30 427
rect -33 389 33 405
rect -33 355 -17 389
rect 17 355 33 389
rect -33 339 33 355
rect -33 281 33 297
rect -33 247 -17 281
rect 17 247 33 281
rect -33 231 33 247
rect -30 209 30 231
rect -30 87 30 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -30 -109 30 -87
rect -30 -231 30 -209
rect -33 -247 33 -231
rect -33 -281 -17 -247
rect 17 -281 33 -247
rect -33 -297 33 -281
rect -33 -355 33 -339
rect -33 -389 -17 -355
rect 17 -389 33 -355
rect -33 -405 33 -389
rect -30 -427 30 -405
rect -30 -549 30 -527
rect -33 -565 33 -549
rect -33 -599 -17 -565
rect 17 -599 33 -565
rect -33 -615 33 -599
<< polycont >>
rect -17 565 17 599
rect -17 355 17 389
rect -17 247 17 281
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -281 17 -247
rect -17 -389 17 -355
rect -17 -599 17 -565
<< locali >>
rect -190 667 -94 701
rect 94 667 190 701
rect -190 605 -156 667
rect 156 605 190 667
rect -33 565 -17 599
rect 17 565 33 599
rect -76 515 -42 531
rect -76 423 -42 439
rect 42 515 76 531
rect 42 423 76 439
rect -33 355 -17 389
rect 17 355 33 389
rect -33 247 -17 281
rect 17 247 33 281
rect -76 197 -42 213
rect -76 105 -42 121
rect 42 197 76 213
rect 42 105 76 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -76 -121 -42 -105
rect -76 -213 -42 -197
rect 42 -121 76 -105
rect 42 -213 76 -197
rect -33 -281 -17 -247
rect 17 -281 33 -247
rect -33 -389 -17 -355
rect 17 -389 33 -355
rect -76 -439 -42 -423
rect -76 -531 -42 -515
rect 42 -439 76 -423
rect 42 -531 76 -515
rect -33 -599 -17 -565
rect 17 -599 33 -565
rect -190 -667 -156 -605
rect 156 -667 190 -605
rect -190 -701 -94 -667
rect 94 -701 190 -667
<< viali >>
rect -17 565 17 599
rect -76 439 -42 515
rect 42 439 76 515
rect -17 355 17 389
rect -17 247 17 281
rect -76 121 -42 197
rect 42 121 76 197
rect -17 37 17 71
rect -17 -71 17 -37
rect -76 -197 -42 -121
rect 42 -197 76 -121
rect -17 -281 17 -247
rect -17 -389 17 -355
rect -76 -515 -42 -439
rect 42 -515 76 -439
rect -17 -599 17 -565
<< metal1 >>
rect -29 599 29 605
rect -29 565 -17 599
rect 17 565 29 599
rect -29 559 29 565
rect -82 515 -36 527
rect -82 439 -76 515
rect -42 439 -36 515
rect -82 427 -36 439
rect 36 515 82 527
rect 36 439 42 515
rect 76 439 82 515
rect 36 427 82 439
rect -29 389 29 395
rect -29 355 -17 389
rect 17 355 29 389
rect -29 349 29 355
rect -29 281 29 287
rect -29 247 -17 281
rect 17 247 29 281
rect -29 241 29 247
rect -82 197 -36 209
rect -82 121 -76 197
rect -42 121 -36 197
rect -82 109 -36 121
rect 36 197 82 209
rect 36 121 42 197
rect 76 121 82 197
rect 36 109 82 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -82 -121 -36 -109
rect -82 -197 -76 -121
rect -42 -197 -36 -121
rect -82 -209 -36 -197
rect 36 -121 82 -109
rect 36 -197 42 -121
rect 76 -197 82 -121
rect 36 -209 82 -197
rect -29 -247 29 -241
rect -29 -281 -17 -247
rect 17 -281 29 -247
rect -29 -287 29 -281
rect -29 -355 29 -349
rect -29 -389 -17 -355
rect 17 -389 29 -355
rect -29 -395 29 -389
rect -82 -439 -36 -427
rect -82 -515 -76 -439
rect -42 -515 -36 -439
rect -82 -527 -36 -515
rect 36 -439 82 -427
rect 36 -515 42 -439
rect 76 -515 82 -439
rect 36 -527 82 -515
rect -29 -565 29 -559
rect -29 -599 -17 -565
rect 17 -599 29 -565
rect -29 -605 29 -599
<< properties >>
string FIXED_BBOX -173 -684 173 684
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.3 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
