magic
tech sky130A
magscale 1 2
timestamp 1729057844
<< error_p >>
rect -29 207 29 213
rect -29 173 -17 207
rect -29 167 29 173
rect -29 -173 29 -167
rect -29 -207 -17 -173
rect -29 -213 29 -207
<< nwell >>
rect -211 -345 211 345
<< pmos >>
rect -15 -126 15 126
<< pdiff >>
rect -73 114 -15 126
rect -73 -114 -61 114
rect -27 -114 -15 114
rect -73 -126 -15 -114
rect 15 114 73 126
rect 15 -114 27 114
rect 61 -114 73 114
rect 15 -126 73 -114
<< pdiffc >>
rect -61 -114 -27 114
rect 27 -114 61 114
<< nsubdiff >>
rect -175 275 -79 309
rect 79 275 175 309
rect -175 213 -141 275
rect 141 213 175 275
rect -175 -275 -141 -213
rect 141 -275 175 -213
rect -175 -309 -79 -275
rect 79 -309 175 -275
<< nsubdiffcont >>
rect -79 275 79 309
rect -175 -213 -141 213
rect 141 -213 175 213
rect -79 -309 79 -275
<< poly >>
rect -33 207 33 223
rect -33 173 -17 207
rect 17 173 33 207
rect -33 157 33 173
rect -15 126 15 157
rect -15 -157 15 -126
rect -33 -173 33 -157
rect -33 -207 -17 -173
rect 17 -207 33 -173
rect -33 -223 33 -207
<< polycont >>
rect -17 173 17 207
rect -17 -207 17 -173
<< locali >>
rect -175 275 -79 309
rect 79 275 175 309
rect -175 213 -141 275
rect 141 213 175 275
rect -33 173 -17 207
rect 17 173 33 207
rect -61 114 -27 130
rect -61 -130 -27 -114
rect 27 114 61 130
rect 27 -130 61 -114
rect -33 -207 -17 -173
rect 17 -207 33 -173
rect -175 -275 -141 -213
rect 141 -275 175 -213
rect -175 -309 -79 -275
rect 79 -309 175 -275
<< viali >>
rect -17 173 17 207
rect -61 -114 -27 114
rect 27 -114 61 114
rect -17 -207 17 -173
<< metal1 >>
rect -29 207 29 213
rect -29 173 -17 207
rect 17 173 29 207
rect -29 167 29 173
rect -67 114 -21 126
rect -67 -114 -61 114
rect -27 -114 -21 114
rect -67 -126 -21 -114
rect 21 114 67 126
rect 21 -114 27 114
rect 61 -114 67 114
rect 21 -126 67 -114
rect -29 -173 29 -167
rect -29 -207 -17 -173
rect 17 -207 29 -173
rect -29 -213 29 -207
<< properties >>
string FIXED_BBOX -158 -292 158 292
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.26 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
