magic
tech sky130A
magscale 1 2
timestamp 1730624594
<< pwell >>
rect -246 -2645 246 2645
<< nmos >>
rect -50 2335 50 2435
rect -50 2017 50 2117
rect -50 1699 50 1799
rect -50 1381 50 1481
rect -50 1063 50 1163
rect -50 745 50 845
rect -50 427 50 527
rect -50 109 50 209
rect -50 -209 50 -109
rect -50 -527 50 -427
rect -50 -845 50 -745
rect -50 -1163 50 -1063
rect -50 -1481 50 -1381
rect -50 -1799 50 -1699
rect -50 -2117 50 -2017
rect -50 -2435 50 -2335
<< ndiff >>
rect -108 2423 -50 2435
rect -108 2347 -96 2423
rect -62 2347 -50 2423
rect -108 2335 -50 2347
rect 50 2423 108 2435
rect 50 2347 62 2423
rect 96 2347 108 2423
rect 50 2335 108 2347
rect -108 2105 -50 2117
rect -108 2029 -96 2105
rect -62 2029 -50 2105
rect -108 2017 -50 2029
rect 50 2105 108 2117
rect 50 2029 62 2105
rect 96 2029 108 2105
rect 50 2017 108 2029
rect -108 1787 -50 1799
rect -108 1711 -96 1787
rect -62 1711 -50 1787
rect -108 1699 -50 1711
rect 50 1787 108 1799
rect 50 1711 62 1787
rect 96 1711 108 1787
rect 50 1699 108 1711
rect -108 1469 -50 1481
rect -108 1393 -96 1469
rect -62 1393 -50 1469
rect -108 1381 -50 1393
rect 50 1469 108 1481
rect 50 1393 62 1469
rect 96 1393 108 1469
rect 50 1381 108 1393
rect -108 1151 -50 1163
rect -108 1075 -96 1151
rect -62 1075 -50 1151
rect -108 1063 -50 1075
rect 50 1151 108 1163
rect 50 1075 62 1151
rect 96 1075 108 1151
rect 50 1063 108 1075
rect -108 833 -50 845
rect -108 757 -96 833
rect -62 757 -50 833
rect -108 745 -50 757
rect 50 833 108 845
rect 50 757 62 833
rect 96 757 108 833
rect 50 745 108 757
rect -108 515 -50 527
rect -108 439 -96 515
rect -62 439 -50 515
rect -108 427 -50 439
rect 50 515 108 527
rect 50 439 62 515
rect 96 439 108 515
rect 50 427 108 439
rect -108 197 -50 209
rect -108 121 -96 197
rect -62 121 -50 197
rect -108 109 -50 121
rect 50 197 108 209
rect 50 121 62 197
rect 96 121 108 197
rect 50 109 108 121
rect -108 -121 -50 -109
rect -108 -197 -96 -121
rect -62 -197 -50 -121
rect -108 -209 -50 -197
rect 50 -121 108 -109
rect 50 -197 62 -121
rect 96 -197 108 -121
rect 50 -209 108 -197
rect -108 -439 -50 -427
rect -108 -515 -96 -439
rect -62 -515 -50 -439
rect -108 -527 -50 -515
rect 50 -439 108 -427
rect 50 -515 62 -439
rect 96 -515 108 -439
rect 50 -527 108 -515
rect -108 -757 -50 -745
rect -108 -833 -96 -757
rect -62 -833 -50 -757
rect -108 -845 -50 -833
rect 50 -757 108 -745
rect 50 -833 62 -757
rect 96 -833 108 -757
rect 50 -845 108 -833
rect -108 -1075 -50 -1063
rect -108 -1151 -96 -1075
rect -62 -1151 -50 -1075
rect -108 -1163 -50 -1151
rect 50 -1075 108 -1063
rect 50 -1151 62 -1075
rect 96 -1151 108 -1075
rect 50 -1163 108 -1151
rect -108 -1393 -50 -1381
rect -108 -1469 -96 -1393
rect -62 -1469 -50 -1393
rect -108 -1481 -50 -1469
rect 50 -1393 108 -1381
rect 50 -1469 62 -1393
rect 96 -1469 108 -1393
rect 50 -1481 108 -1469
rect -108 -1711 -50 -1699
rect -108 -1787 -96 -1711
rect -62 -1787 -50 -1711
rect -108 -1799 -50 -1787
rect 50 -1711 108 -1699
rect 50 -1787 62 -1711
rect 96 -1787 108 -1711
rect 50 -1799 108 -1787
rect -108 -2029 -50 -2017
rect -108 -2105 -96 -2029
rect -62 -2105 -50 -2029
rect -108 -2117 -50 -2105
rect 50 -2029 108 -2017
rect 50 -2105 62 -2029
rect 96 -2105 108 -2029
rect 50 -2117 108 -2105
rect -108 -2347 -50 -2335
rect -108 -2423 -96 -2347
rect -62 -2423 -50 -2347
rect -108 -2435 -50 -2423
rect 50 -2347 108 -2335
rect 50 -2423 62 -2347
rect 96 -2423 108 -2347
rect 50 -2435 108 -2423
<< ndiffc >>
rect -96 2347 -62 2423
rect 62 2347 96 2423
rect -96 2029 -62 2105
rect 62 2029 96 2105
rect -96 1711 -62 1787
rect 62 1711 96 1787
rect -96 1393 -62 1469
rect 62 1393 96 1469
rect -96 1075 -62 1151
rect 62 1075 96 1151
rect -96 757 -62 833
rect 62 757 96 833
rect -96 439 -62 515
rect 62 439 96 515
rect -96 121 -62 197
rect 62 121 96 197
rect -96 -197 -62 -121
rect 62 -197 96 -121
rect -96 -515 -62 -439
rect 62 -515 96 -439
rect -96 -833 -62 -757
rect 62 -833 96 -757
rect -96 -1151 -62 -1075
rect 62 -1151 96 -1075
rect -96 -1469 -62 -1393
rect 62 -1469 96 -1393
rect -96 -1787 -62 -1711
rect 62 -1787 96 -1711
rect -96 -2105 -62 -2029
rect 62 -2105 96 -2029
rect -96 -2423 -62 -2347
rect 62 -2423 96 -2347
<< psubdiff >>
rect -210 2575 -114 2609
rect 114 2575 210 2609
rect -210 2513 -176 2575
rect 176 2513 210 2575
rect -210 -2575 -176 -2513
rect 176 -2575 210 -2513
rect -210 -2609 -114 -2575
rect 114 -2609 210 -2575
<< psubdiffcont >>
rect -114 2575 114 2609
rect -210 -2513 -176 2513
rect 176 -2513 210 2513
rect -114 -2609 114 -2575
<< poly >>
rect -50 2507 50 2523
rect -50 2473 -34 2507
rect 34 2473 50 2507
rect -50 2435 50 2473
rect -50 2297 50 2335
rect -50 2263 -34 2297
rect 34 2263 50 2297
rect -50 2247 50 2263
rect -50 2189 50 2205
rect -50 2155 -34 2189
rect 34 2155 50 2189
rect -50 2117 50 2155
rect -50 1979 50 2017
rect -50 1945 -34 1979
rect 34 1945 50 1979
rect -50 1929 50 1945
rect -50 1871 50 1887
rect -50 1837 -34 1871
rect 34 1837 50 1871
rect -50 1799 50 1837
rect -50 1661 50 1699
rect -50 1627 -34 1661
rect 34 1627 50 1661
rect -50 1611 50 1627
rect -50 1553 50 1569
rect -50 1519 -34 1553
rect 34 1519 50 1553
rect -50 1481 50 1519
rect -50 1343 50 1381
rect -50 1309 -34 1343
rect 34 1309 50 1343
rect -50 1293 50 1309
rect -50 1235 50 1251
rect -50 1201 -34 1235
rect 34 1201 50 1235
rect -50 1163 50 1201
rect -50 1025 50 1063
rect -50 991 -34 1025
rect 34 991 50 1025
rect -50 975 50 991
rect -50 917 50 933
rect -50 883 -34 917
rect 34 883 50 917
rect -50 845 50 883
rect -50 707 50 745
rect -50 673 -34 707
rect 34 673 50 707
rect -50 657 50 673
rect -50 599 50 615
rect -50 565 -34 599
rect 34 565 50 599
rect -50 527 50 565
rect -50 389 50 427
rect -50 355 -34 389
rect 34 355 50 389
rect -50 339 50 355
rect -50 281 50 297
rect -50 247 -34 281
rect 34 247 50 281
rect -50 209 50 247
rect -50 71 50 109
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -109 50 -71
rect -50 -247 50 -209
rect -50 -281 -34 -247
rect 34 -281 50 -247
rect -50 -297 50 -281
rect -50 -355 50 -339
rect -50 -389 -34 -355
rect 34 -389 50 -355
rect -50 -427 50 -389
rect -50 -565 50 -527
rect -50 -599 -34 -565
rect 34 -599 50 -565
rect -50 -615 50 -599
rect -50 -673 50 -657
rect -50 -707 -34 -673
rect 34 -707 50 -673
rect -50 -745 50 -707
rect -50 -883 50 -845
rect -50 -917 -34 -883
rect 34 -917 50 -883
rect -50 -933 50 -917
rect -50 -991 50 -975
rect -50 -1025 -34 -991
rect 34 -1025 50 -991
rect -50 -1063 50 -1025
rect -50 -1201 50 -1163
rect -50 -1235 -34 -1201
rect 34 -1235 50 -1201
rect -50 -1251 50 -1235
rect -50 -1309 50 -1293
rect -50 -1343 -34 -1309
rect 34 -1343 50 -1309
rect -50 -1381 50 -1343
rect -50 -1519 50 -1481
rect -50 -1553 -34 -1519
rect 34 -1553 50 -1519
rect -50 -1569 50 -1553
rect -50 -1627 50 -1611
rect -50 -1661 -34 -1627
rect 34 -1661 50 -1627
rect -50 -1699 50 -1661
rect -50 -1837 50 -1799
rect -50 -1871 -34 -1837
rect 34 -1871 50 -1837
rect -50 -1887 50 -1871
rect -50 -1945 50 -1929
rect -50 -1979 -34 -1945
rect 34 -1979 50 -1945
rect -50 -2017 50 -1979
rect -50 -2155 50 -2117
rect -50 -2189 -34 -2155
rect 34 -2189 50 -2155
rect -50 -2205 50 -2189
rect -50 -2263 50 -2247
rect -50 -2297 -34 -2263
rect 34 -2297 50 -2263
rect -50 -2335 50 -2297
rect -50 -2473 50 -2435
rect -50 -2507 -34 -2473
rect 34 -2507 50 -2473
rect -50 -2523 50 -2507
<< polycont >>
rect -34 2473 34 2507
rect -34 2263 34 2297
rect -34 2155 34 2189
rect -34 1945 34 1979
rect -34 1837 34 1871
rect -34 1627 34 1661
rect -34 1519 34 1553
rect -34 1309 34 1343
rect -34 1201 34 1235
rect -34 991 34 1025
rect -34 883 34 917
rect -34 673 34 707
rect -34 565 34 599
rect -34 355 34 389
rect -34 247 34 281
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -281 34 -247
rect -34 -389 34 -355
rect -34 -599 34 -565
rect -34 -707 34 -673
rect -34 -917 34 -883
rect -34 -1025 34 -991
rect -34 -1235 34 -1201
rect -34 -1343 34 -1309
rect -34 -1553 34 -1519
rect -34 -1661 34 -1627
rect -34 -1871 34 -1837
rect -34 -1979 34 -1945
rect -34 -2189 34 -2155
rect -34 -2297 34 -2263
rect -34 -2507 34 -2473
<< locali >>
rect -210 2575 -114 2609
rect 114 2575 210 2609
rect -210 2513 -176 2575
rect 176 2513 210 2575
rect -50 2473 -34 2507
rect 34 2473 50 2507
rect -96 2423 -62 2439
rect -96 2331 -62 2347
rect 62 2423 96 2439
rect 62 2331 96 2347
rect -50 2263 -34 2297
rect 34 2263 50 2297
rect -50 2155 -34 2189
rect 34 2155 50 2189
rect -96 2105 -62 2121
rect -96 2013 -62 2029
rect 62 2105 96 2121
rect 62 2013 96 2029
rect -50 1945 -34 1979
rect 34 1945 50 1979
rect -50 1837 -34 1871
rect 34 1837 50 1871
rect -96 1787 -62 1803
rect -96 1695 -62 1711
rect 62 1787 96 1803
rect 62 1695 96 1711
rect -50 1627 -34 1661
rect 34 1627 50 1661
rect -50 1519 -34 1553
rect 34 1519 50 1553
rect -96 1469 -62 1485
rect -96 1377 -62 1393
rect 62 1469 96 1485
rect 62 1377 96 1393
rect -50 1309 -34 1343
rect 34 1309 50 1343
rect -50 1201 -34 1235
rect 34 1201 50 1235
rect -96 1151 -62 1167
rect -96 1059 -62 1075
rect 62 1151 96 1167
rect 62 1059 96 1075
rect -50 991 -34 1025
rect 34 991 50 1025
rect -50 883 -34 917
rect 34 883 50 917
rect -96 833 -62 849
rect -96 741 -62 757
rect 62 833 96 849
rect 62 741 96 757
rect -50 673 -34 707
rect 34 673 50 707
rect -50 565 -34 599
rect 34 565 50 599
rect -96 515 -62 531
rect -96 423 -62 439
rect 62 515 96 531
rect 62 423 96 439
rect -50 355 -34 389
rect 34 355 50 389
rect -50 247 -34 281
rect 34 247 50 281
rect -96 197 -62 213
rect -96 105 -62 121
rect 62 197 96 213
rect 62 105 96 121
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -121 -62 -105
rect -96 -213 -62 -197
rect 62 -121 96 -105
rect 62 -213 96 -197
rect -50 -281 -34 -247
rect 34 -281 50 -247
rect -50 -389 -34 -355
rect 34 -389 50 -355
rect -96 -439 -62 -423
rect -96 -531 -62 -515
rect 62 -439 96 -423
rect 62 -531 96 -515
rect -50 -599 -34 -565
rect 34 -599 50 -565
rect -50 -707 -34 -673
rect 34 -707 50 -673
rect -96 -757 -62 -741
rect -96 -849 -62 -833
rect 62 -757 96 -741
rect 62 -849 96 -833
rect -50 -917 -34 -883
rect 34 -917 50 -883
rect -50 -1025 -34 -991
rect 34 -1025 50 -991
rect -96 -1075 -62 -1059
rect -96 -1167 -62 -1151
rect 62 -1075 96 -1059
rect 62 -1167 96 -1151
rect -50 -1235 -34 -1201
rect 34 -1235 50 -1201
rect -50 -1343 -34 -1309
rect 34 -1343 50 -1309
rect -96 -1393 -62 -1377
rect -96 -1485 -62 -1469
rect 62 -1393 96 -1377
rect 62 -1485 96 -1469
rect -50 -1553 -34 -1519
rect 34 -1553 50 -1519
rect -50 -1661 -34 -1627
rect 34 -1661 50 -1627
rect -96 -1711 -62 -1695
rect -96 -1803 -62 -1787
rect 62 -1711 96 -1695
rect 62 -1803 96 -1787
rect -50 -1871 -34 -1837
rect 34 -1871 50 -1837
rect -50 -1979 -34 -1945
rect 34 -1979 50 -1945
rect -96 -2029 -62 -2013
rect -96 -2121 -62 -2105
rect 62 -2029 96 -2013
rect 62 -2121 96 -2105
rect -50 -2189 -34 -2155
rect 34 -2189 50 -2155
rect -50 -2297 -34 -2263
rect 34 -2297 50 -2263
rect -96 -2347 -62 -2331
rect -96 -2439 -62 -2423
rect 62 -2347 96 -2331
rect 62 -2439 96 -2423
rect -50 -2507 -34 -2473
rect 34 -2507 50 -2473
rect -210 -2575 -176 -2513
rect 176 -2575 210 -2513
rect -210 -2609 -114 -2575
rect 114 -2609 210 -2575
<< viali >>
rect -34 2473 34 2507
rect -96 2347 -62 2423
rect 62 2347 96 2423
rect -34 2263 34 2297
rect -34 2155 34 2189
rect -96 2029 -62 2105
rect 62 2029 96 2105
rect -34 1945 34 1979
rect -34 1837 34 1871
rect -96 1711 -62 1787
rect 62 1711 96 1787
rect -34 1627 34 1661
rect -34 1519 34 1553
rect -96 1393 -62 1469
rect 62 1393 96 1469
rect -34 1309 34 1343
rect -34 1201 34 1235
rect -96 1075 -62 1151
rect 62 1075 96 1151
rect -34 991 34 1025
rect -34 883 34 917
rect -96 757 -62 833
rect 62 757 96 833
rect -34 673 34 707
rect -34 565 34 599
rect -96 439 -62 515
rect 62 439 96 515
rect -34 355 34 389
rect -34 247 34 281
rect -96 121 -62 197
rect 62 121 96 197
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -197 -62 -121
rect 62 -197 96 -121
rect -34 -281 34 -247
rect -34 -389 34 -355
rect -96 -515 -62 -439
rect 62 -515 96 -439
rect -34 -599 34 -565
rect -34 -707 34 -673
rect -96 -833 -62 -757
rect 62 -833 96 -757
rect -34 -917 34 -883
rect -34 -1025 34 -991
rect -96 -1151 -62 -1075
rect 62 -1151 96 -1075
rect -34 -1235 34 -1201
rect -34 -1343 34 -1309
rect -96 -1469 -62 -1393
rect 62 -1469 96 -1393
rect -34 -1553 34 -1519
rect -34 -1661 34 -1627
rect -96 -1787 -62 -1711
rect 62 -1787 96 -1711
rect -34 -1871 34 -1837
rect -34 -1979 34 -1945
rect -96 -2105 -62 -2029
rect 62 -2105 96 -2029
rect -34 -2189 34 -2155
rect -34 -2297 34 -2263
rect -96 -2423 -62 -2347
rect 62 -2423 96 -2347
rect -34 -2507 34 -2473
<< metal1 >>
rect -46 2507 46 2513
rect -46 2473 -34 2507
rect 34 2473 46 2507
rect -46 2467 46 2473
rect -102 2423 -56 2435
rect -102 2347 -96 2423
rect -62 2347 -56 2423
rect -102 2335 -56 2347
rect 56 2423 102 2435
rect 56 2347 62 2423
rect 96 2347 102 2423
rect 56 2335 102 2347
rect -46 2297 46 2303
rect -46 2263 -34 2297
rect 34 2263 46 2297
rect -46 2257 46 2263
rect -46 2189 46 2195
rect -46 2155 -34 2189
rect 34 2155 46 2189
rect -46 2149 46 2155
rect -102 2105 -56 2117
rect -102 2029 -96 2105
rect -62 2029 -56 2105
rect -102 2017 -56 2029
rect 56 2105 102 2117
rect 56 2029 62 2105
rect 96 2029 102 2105
rect 56 2017 102 2029
rect -46 1979 46 1985
rect -46 1945 -34 1979
rect 34 1945 46 1979
rect -46 1939 46 1945
rect -46 1871 46 1877
rect -46 1837 -34 1871
rect 34 1837 46 1871
rect -46 1831 46 1837
rect -102 1787 -56 1799
rect -102 1711 -96 1787
rect -62 1711 -56 1787
rect -102 1699 -56 1711
rect 56 1787 102 1799
rect 56 1711 62 1787
rect 96 1711 102 1787
rect 56 1699 102 1711
rect -46 1661 46 1667
rect -46 1627 -34 1661
rect 34 1627 46 1661
rect -46 1621 46 1627
rect -46 1553 46 1559
rect -46 1519 -34 1553
rect 34 1519 46 1553
rect -46 1513 46 1519
rect -102 1469 -56 1481
rect -102 1393 -96 1469
rect -62 1393 -56 1469
rect -102 1381 -56 1393
rect 56 1469 102 1481
rect 56 1393 62 1469
rect 96 1393 102 1469
rect 56 1381 102 1393
rect -46 1343 46 1349
rect -46 1309 -34 1343
rect 34 1309 46 1343
rect -46 1303 46 1309
rect -46 1235 46 1241
rect -46 1201 -34 1235
rect 34 1201 46 1235
rect -46 1195 46 1201
rect -102 1151 -56 1163
rect -102 1075 -96 1151
rect -62 1075 -56 1151
rect -102 1063 -56 1075
rect 56 1151 102 1163
rect 56 1075 62 1151
rect 96 1075 102 1151
rect 56 1063 102 1075
rect -46 1025 46 1031
rect -46 991 -34 1025
rect 34 991 46 1025
rect -46 985 46 991
rect -46 917 46 923
rect -46 883 -34 917
rect 34 883 46 917
rect -46 877 46 883
rect -102 833 -56 845
rect -102 757 -96 833
rect -62 757 -56 833
rect -102 745 -56 757
rect 56 833 102 845
rect 56 757 62 833
rect 96 757 102 833
rect 56 745 102 757
rect -46 707 46 713
rect -46 673 -34 707
rect 34 673 46 707
rect -46 667 46 673
rect -46 599 46 605
rect -46 565 -34 599
rect 34 565 46 599
rect -46 559 46 565
rect -102 515 -56 527
rect -102 439 -96 515
rect -62 439 -56 515
rect -102 427 -56 439
rect 56 515 102 527
rect 56 439 62 515
rect 96 439 102 515
rect 56 427 102 439
rect -46 389 46 395
rect -46 355 -34 389
rect 34 355 46 389
rect -46 349 46 355
rect -46 281 46 287
rect -46 247 -34 281
rect 34 247 46 281
rect -46 241 46 247
rect -102 197 -56 209
rect -102 121 -96 197
rect -62 121 -56 197
rect -102 109 -56 121
rect 56 197 102 209
rect 56 121 62 197
rect 96 121 102 197
rect 56 109 102 121
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -121 -56 -109
rect -102 -197 -96 -121
rect -62 -197 -56 -121
rect -102 -209 -56 -197
rect 56 -121 102 -109
rect 56 -197 62 -121
rect 96 -197 102 -121
rect 56 -209 102 -197
rect -46 -247 46 -241
rect -46 -281 -34 -247
rect 34 -281 46 -247
rect -46 -287 46 -281
rect -46 -355 46 -349
rect -46 -389 -34 -355
rect 34 -389 46 -355
rect -46 -395 46 -389
rect -102 -439 -56 -427
rect -102 -515 -96 -439
rect -62 -515 -56 -439
rect -102 -527 -56 -515
rect 56 -439 102 -427
rect 56 -515 62 -439
rect 96 -515 102 -439
rect 56 -527 102 -515
rect -46 -565 46 -559
rect -46 -599 -34 -565
rect 34 -599 46 -565
rect -46 -605 46 -599
rect -46 -673 46 -667
rect -46 -707 -34 -673
rect 34 -707 46 -673
rect -46 -713 46 -707
rect -102 -757 -56 -745
rect -102 -833 -96 -757
rect -62 -833 -56 -757
rect -102 -845 -56 -833
rect 56 -757 102 -745
rect 56 -833 62 -757
rect 96 -833 102 -757
rect 56 -845 102 -833
rect -46 -883 46 -877
rect -46 -917 -34 -883
rect 34 -917 46 -883
rect -46 -923 46 -917
rect -46 -991 46 -985
rect -46 -1025 -34 -991
rect 34 -1025 46 -991
rect -46 -1031 46 -1025
rect -102 -1075 -56 -1063
rect -102 -1151 -96 -1075
rect -62 -1151 -56 -1075
rect -102 -1163 -56 -1151
rect 56 -1075 102 -1063
rect 56 -1151 62 -1075
rect 96 -1151 102 -1075
rect 56 -1163 102 -1151
rect -46 -1201 46 -1195
rect -46 -1235 -34 -1201
rect 34 -1235 46 -1201
rect -46 -1241 46 -1235
rect -46 -1309 46 -1303
rect -46 -1343 -34 -1309
rect 34 -1343 46 -1309
rect -46 -1349 46 -1343
rect -102 -1393 -56 -1381
rect -102 -1469 -96 -1393
rect -62 -1469 -56 -1393
rect -102 -1481 -56 -1469
rect 56 -1393 102 -1381
rect 56 -1469 62 -1393
rect 96 -1469 102 -1393
rect 56 -1481 102 -1469
rect -46 -1519 46 -1513
rect -46 -1553 -34 -1519
rect 34 -1553 46 -1519
rect -46 -1559 46 -1553
rect -46 -1627 46 -1621
rect -46 -1661 -34 -1627
rect 34 -1661 46 -1627
rect -46 -1667 46 -1661
rect -102 -1711 -56 -1699
rect -102 -1787 -96 -1711
rect -62 -1787 -56 -1711
rect -102 -1799 -56 -1787
rect 56 -1711 102 -1699
rect 56 -1787 62 -1711
rect 96 -1787 102 -1711
rect 56 -1799 102 -1787
rect -46 -1837 46 -1831
rect -46 -1871 -34 -1837
rect 34 -1871 46 -1837
rect -46 -1877 46 -1871
rect -46 -1945 46 -1939
rect -46 -1979 -34 -1945
rect 34 -1979 46 -1945
rect -46 -1985 46 -1979
rect -102 -2029 -56 -2017
rect -102 -2105 -96 -2029
rect -62 -2105 -56 -2029
rect -102 -2117 -56 -2105
rect 56 -2029 102 -2017
rect 56 -2105 62 -2029
rect 96 -2105 102 -2029
rect 56 -2117 102 -2105
rect -46 -2155 46 -2149
rect -46 -2189 -34 -2155
rect 34 -2189 46 -2155
rect -46 -2195 46 -2189
rect -46 -2263 46 -2257
rect -46 -2297 -34 -2263
rect 34 -2297 46 -2263
rect -46 -2303 46 -2297
rect -102 -2347 -56 -2335
rect -102 -2423 -96 -2347
rect -62 -2423 -56 -2347
rect -102 -2435 -56 -2423
rect 56 -2347 102 -2335
rect 56 -2423 62 -2347
rect 96 -2423 102 -2347
rect 56 -2435 102 -2423
rect -46 -2473 46 -2467
rect -46 -2507 -34 -2473
rect 34 -2507 46 -2473
rect -46 -2513 46 -2507
<< properties >>
string FIXED_BBOX -193 -2592 193 2592
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.5 m 16 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
