magic
tech sky130A
magscale 1 2
timestamp 1731265361
<< locali >>
rect -106 1173 9858 1175
rect -106 1139 61 1173
rect 95 1139 133 1173
rect 167 1139 205 1173
rect 239 1139 277 1173
rect 311 1139 349 1173
rect 383 1139 421 1173
rect 455 1139 493 1173
rect 527 1139 565 1173
rect 599 1139 637 1173
rect 671 1139 709 1173
rect 743 1139 781 1173
rect 815 1139 853 1173
rect 887 1139 925 1173
rect 959 1139 997 1173
rect 1031 1139 1069 1173
rect 1103 1139 1141 1173
rect 1175 1139 1213 1173
rect 1247 1139 1285 1173
rect 1319 1139 1357 1173
rect 1391 1139 1429 1173
rect 1463 1139 1501 1173
rect 1535 1139 1573 1173
rect 1607 1139 1645 1173
rect 1679 1139 1717 1173
rect 1751 1139 1789 1173
rect 1823 1139 1861 1173
rect 1895 1139 1933 1173
rect 1967 1139 2005 1173
rect 2039 1139 2077 1173
rect 2111 1139 2149 1173
rect 2183 1139 2221 1173
rect 2255 1139 2293 1173
rect 2327 1139 2365 1173
rect 2399 1139 2437 1173
rect 2471 1139 2509 1173
rect 2543 1139 2581 1173
rect 2615 1139 2653 1173
rect 2687 1139 2725 1173
rect 2759 1139 2797 1173
rect 2831 1139 2869 1173
rect 2903 1139 2941 1173
rect 2975 1139 3013 1173
rect 3047 1139 3085 1173
rect 3119 1139 3347 1173
rect 3381 1139 3419 1173
rect 3453 1139 3491 1173
rect 3525 1139 3563 1173
rect 3597 1139 3635 1173
rect 3669 1139 3707 1173
rect 3741 1139 3779 1173
rect 3813 1139 3851 1173
rect 3885 1139 3923 1173
rect 3957 1139 3995 1173
rect 4029 1139 4067 1173
rect 4101 1139 4139 1173
rect 4173 1139 4211 1173
rect 4245 1139 4283 1173
rect 4317 1139 4355 1173
rect 4389 1139 4427 1173
rect 4461 1139 4499 1173
rect 4533 1139 4571 1173
rect 4605 1139 4643 1173
rect 4677 1139 4715 1173
rect 4749 1139 4787 1173
rect 4821 1139 4859 1173
rect 4893 1139 4931 1173
rect 4965 1139 5003 1173
rect 5037 1139 5075 1173
rect 5109 1139 5147 1173
rect 5181 1139 5219 1173
rect 5253 1139 5291 1173
rect 5325 1139 5363 1173
rect 5397 1139 5435 1173
rect 5469 1139 5507 1173
rect 5541 1139 5579 1173
rect 5613 1139 5651 1173
rect 5685 1139 5723 1173
rect 5757 1139 5795 1173
rect 5829 1139 5867 1173
rect 5901 1139 5939 1173
rect 5973 1139 6011 1173
rect 6045 1139 6083 1173
rect 6117 1139 6155 1173
rect 6189 1139 6227 1173
rect 6261 1139 6299 1173
rect 6333 1139 6371 1173
rect 6405 1139 6633 1173
rect 6667 1139 6705 1173
rect 6739 1139 6777 1173
rect 6811 1139 6849 1173
rect 6883 1139 6921 1173
rect 6955 1139 6993 1173
rect 7027 1139 7065 1173
rect 7099 1139 7137 1173
rect 7171 1139 7209 1173
rect 7243 1139 7281 1173
rect 7315 1139 7353 1173
rect 7387 1139 7425 1173
rect 7459 1139 7497 1173
rect 7531 1139 7569 1173
rect 7603 1139 7641 1173
rect 7675 1139 7713 1173
rect 7747 1139 7785 1173
rect 7819 1139 7857 1173
rect 7891 1139 7929 1173
rect 7963 1139 8001 1173
rect 8035 1139 8073 1173
rect 8107 1139 8145 1173
rect 8179 1139 8217 1173
rect 8251 1139 8289 1173
rect 8323 1139 8361 1173
rect 8395 1139 8433 1173
rect 8467 1139 8505 1173
rect 8539 1139 8577 1173
rect 8611 1139 8649 1173
rect 8683 1139 8721 1173
rect 8755 1139 8793 1173
rect 8827 1139 8865 1173
rect 8899 1139 8937 1173
rect 8971 1139 9009 1173
rect 9043 1139 9081 1173
rect 9115 1139 9153 1173
rect 9187 1139 9225 1173
rect 9259 1139 9297 1173
rect 9331 1139 9369 1173
rect 9403 1139 9441 1173
rect 9475 1139 9513 1173
rect 9547 1139 9585 1173
rect 9619 1139 9657 1173
rect 9691 1139 9858 1173
rect -106 1105 9858 1139
rect -106 -427 -36 1105
rect 6502 1021 6536 1043
rect 6502 949 6536 987
rect 6502 877 6536 915
rect 6502 805 6536 843
rect 6502 733 6536 771
rect 6502 661 6536 699
rect 6502 589 6536 627
rect 6502 517 6536 555
rect 6502 445 6536 483
rect 6502 373 6536 411
rect 6502 301 6536 339
rect 6502 229 6536 267
rect 6502 157 6536 195
rect 6502 85 6536 123
rect 6502 13 6536 51
rect 6502 -59 6536 -21
rect 6502 -131 6536 -93
rect 6502 -203 6536 -165
rect 6502 -275 6536 -237
rect 6502 -331 6536 -309
rect 9788 -427 9858 1105
rect -107 -1577 -37 -863
rect 9787 -1577 9857 -863
rect -107 -1647 9857 -1577
rect -107 -1680 9893 -1647
rect -107 -1714 -92 -1680
rect -58 -1714 -20 -1680
rect 14 -1714 52 -1680
rect 86 -1714 124 -1680
rect 158 -1714 196 -1680
rect 230 -1714 268 -1680
rect 302 -1714 340 -1680
rect 374 -1714 412 -1680
rect 446 -1714 484 -1680
rect 518 -1714 556 -1680
rect 590 -1714 628 -1680
rect 662 -1714 700 -1680
rect 734 -1714 772 -1680
rect 806 -1714 844 -1680
rect 878 -1714 916 -1680
rect 950 -1714 988 -1680
rect 1022 -1714 1060 -1680
rect 1094 -1714 1132 -1680
rect 1166 -1714 1204 -1680
rect 1238 -1714 1276 -1680
rect 1310 -1714 1348 -1680
rect 1382 -1714 1420 -1680
rect 1454 -1714 1492 -1680
rect 1526 -1714 1564 -1680
rect 1598 -1714 1636 -1680
rect 1670 -1714 1708 -1680
rect 1742 -1714 1780 -1680
rect 1814 -1714 1852 -1680
rect 1886 -1714 1924 -1680
rect 1958 -1714 1996 -1680
rect 2030 -1714 2068 -1680
rect 2102 -1714 2140 -1680
rect 2174 -1714 2212 -1680
rect 2246 -1714 2284 -1680
rect 2318 -1714 2356 -1680
rect 2390 -1714 2428 -1680
rect 2462 -1714 2500 -1680
rect 2534 -1714 2572 -1680
rect 2606 -1714 2644 -1680
rect 2678 -1714 2716 -1680
rect 2750 -1714 2788 -1680
rect 2822 -1714 2860 -1680
rect 2894 -1714 2932 -1680
rect 2966 -1714 3004 -1680
rect 3038 -1714 3076 -1680
rect 3110 -1714 3148 -1680
rect 3182 -1714 3220 -1680
rect 3254 -1714 3292 -1680
rect 3326 -1714 3364 -1680
rect 3398 -1714 3436 -1680
rect 3470 -1714 3508 -1680
rect 3542 -1714 3580 -1680
rect 3614 -1714 3652 -1680
rect 3686 -1714 3724 -1680
rect 3758 -1714 3796 -1680
rect 3830 -1714 3868 -1680
rect 3902 -1714 3940 -1680
rect 3974 -1714 4012 -1680
rect 4046 -1714 4084 -1680
rect 4118 -1714 4156 -1680
rect 4190 -1714 4228 -1680
rect 4262 -1714 4300 -1680
rect 4334 -1714 4372 -1680
rect 4406 -1714 4444 -1680
rect 4478 -1714 4516 -1680
rect 4550 -1714 4588 -1680
rect 4622 -1714 4660 -1680
rect 4694 -1714 4732 -1680
rect 4766 -1714 4804 -1680
rect 4838 -1714 4876 -1680
rect 4910 -1714 4948 -1680
rect 4982 -1714 5020 -1680
rect 5054 -1714 5092 -1680
rect 5126 -1714 5164 -1680
rect 5198 -1714 5236 -1680
rect 5270 -1714 5308 -1680
rect 5342 -1714 5380 -1680
rect 5414 -1714 5452 -1680
rect 5486 -1714 5524 -1680
rect 5558 -1714 5596 -1680
rect 5630 -1714 5668 -1680
rect 5702 -1714 5740 -1680
rect 5774 -1714 5812 -1680
rect 5846 -1714 5884 -1680
rect 5918 -1714 5956 -1680
rect 5990 -1714 6028 -1680
rect 6062 -1714 6100 -1680
rect 6134 -1714 6172 -1680
rect 6206 -1714 6244 -1680
rect 6278 -1714 6316 -1680
rect 6350 -1714 6388 -1680
rect 6422 -1714 6460 -1680
rect 6494 -1714 6532 -1680
rect 6566 -1714 6604 -1680
rect 6638 -1714 6676 -1680
rect 6710 -1714 6748 -1680
rect 6782 -1714 6820 -1680
rect 6854 -1714 6892 -1680
rect 6926 -1714 6964 -1680
rect 6998 -1714 7036 -1680
rect 7070 -1714 7108 -1680
rect 7142 -1714 7180 -1680
rect 7214 -1714 7252 -1680
rect 7286 -1714 7324 -1680
rect 7358 -1714 7396 -1680
rect 7430 -1714 7468 -1680
rect 7502 -1714 7540 -1680
rect 7574 -1714 7612 -1680
rect 7646 -1714 7684 -1680
rect 7718 -1714 7756 -1680
rect 7790 -1714 7828 -1680
rect 7862 -1714 7900 -1680
rect 7934 -1714 7972 -1680
rect 8006 -1714 8044 -1680
rect 8078 -1714 8116 -1680
rect 8150 -1714 8188 -1680
rect 8222 -1714 8260 -1680
rect 8294 -1714 8332 -1680
rect 8366 -1714 8404 -1680
rect 8438 -1714 8476 -1680
rect 8510 -1714 8548 -1680
rect 8582 -1714 8620 -1680
rect 8654 -1714 8692 -1680
rect 8726 -1714 8764 -1680
rect 8798 -1714 8836 -1680
rect 8870 -1714 8908 -1680
rect 8942 -1714 8980 -1680
rect 9014 -1714 9052 -1680
rect 9086 -1714 9124 -1680
rect 9158 -1714 9196 -1680
rect 9230 -1714 9268 -1680
rect 9302 -1714 9340 -1680
rect 9374 -1714 9412 -1680
rect 9446 -1714 9484 -1680
rect 9518 -1714 9556 -1680
rect 9590 -1714 9628 -1680
rect 9662 -1714 9700 -1680
rect 9734 -1714 9772 -1680
rect 9806 -1714 9844 -1680
rect 9878 -1714 9893 -1680
rect -107 -1747 9893 -1714
<< viali >>
rect 61 1139 95 1173
rect 133 1139 167 1173
rect 205 1139 239 1173
rect 277 1139 311 1173
rect 349 1139 383 1173
rect 421 1139 455 1173
rect 493 1139 527 1173
rect 565 1139 599 1173
rect 637 1139 671 1173
rect 709 1139 743 1173
rect 781 1139 815 1173
rect 853 1139 887 1173
rect 925 1139 959 1173
rect 997 1139 1031 1173
rect 1069 1139 1103 1173
rect 1141 1139 1175 1173
rect 1213 1139 1247 1173
rect 1285 1139 1319 1173
rect 1357 1139 1391 1173
rect 1429 1139 1463 1173
rect 1501 1139 1535 1173
rect 1573 1139 1607 1173
rect 1645 1139 1679 1173
rect 1717 1139 1751 1173
rect 1789 1139 1823 1173
rect 1861 1139 1895 1173
rect 1933 1139 1967 1173
rect 2005 1139 2039 1173
rect 2077 1139 2111 1173
rect 2149 1139 2183 1173
rect 2221 1139 2255 1173
rect 2293 1139 2327 1173
rect 2365 1139 2399 1173
rect 2437 1139 2471 1173
rect 2509 1139 2543 1173
rect 2581 1139 2615 1173
rect 2653 1139 2687 1173
rect 2725 1139 2759 1173
rect 2797 1139 2831 1173
rect 2869 1139 2903 1173
rect 2941 1139 2975 1173
rect 3013 1139 3047 1173
rect 3085 1139 3119 1173
rect 3347 1139 3381 1173
rect 3419 1139 3453 1173
rect 3491 1139 3525 1173
rect 3563 1139 3597 1173
rect 3635 1139 3669 1173
rect 3707 1139 3741 1173
rect 3779 1139 3813 1173
rect 3851 1139 3885 1173
rect 3923 1139 3957 1173
rect 3995 1139 4029 1173
rect 4067 1139 4101 1173
rect 4139 1139 4173 1173
rect 4211 1139 4245 1173
rect 4283 1139 4317 1173
rect 4355 1139 4389 1173
rect 4427 1139 4461 1173
rect 4499 1139 4533 1173
rect 4571 1139 4605 1173
rect 4643 1139 4677 1173
rect 4715 1139 4749 1173
rect 4787 1139 4821 1173
rect 4859 1139 4893 1173
rect 4931 1139 4965 1173
rect 5003 1139 5037 1173
rect 5075 1139 5109 1173
rect 5147 1139 5181 1173
rect 5219 1139 5253 1173
rect 5291 1139 5325 1173
rect 5363 1139 5397 1173
rect 5435 1139 5469 1173
rect 5507 1139 5541 1173
rect 5579 1139 5613 1173
rect 5651 1139 5685 1173
rect 5723 1139 5757 1173
rect 5795 1139 5829 1173
rect 5867 1139 5901 1173
rect 5939 1139 5973 1173
rect 6011 1139 6045 1173
rect 6083 1139 6117 1173
rect 6155 1139 6189 1173
rect 6227 1139 6261 1173
rect 6299 1139 6333 1173
rect 6371 1139 6405 1173
rect 6633 1139 6667 1173
rect 6705 1139 6739 1173
rect 6777 1139 6811 1173
rect 6849 1139 6883 1173
rect 6921 1139 6955 1173
rect 6993 1139 7027 1173
rect 7065 1139 7099 1173
rect 7137 1139 7171 1173
rect 7209 1139 7243 1173
rect 7281 1139 7315 1173
rect 7353 1139 7387 1173
rect 7425 1139 7459 1173
rect 7497 1139 7531 1173
rect 7569 1139 7603 1173
rect 7641 1139 7675 1173
rect 7713 1139 7747 1173
rect 7785 1139 7819 1173
rect 7857 1139 7891 1173
rect 7929 1139 7963 1173
rect 8001 1139 8035 1173
rect 8073 1139 8107 1173
rect 8145 1139 8179 1173
rect 8217 1139 8251 1173
rect 8289 1139 8323 1173
rect 8361 1139 8395 1173
rect 8433 1139 8467 1173
rect 8505 1139 8539 1173
rect 8577 1139 8611 1173
rect 8649 1139 8683 1173
rect 8721 1139 8755 1173
rect 8793 1139 8827 1173
rect 8865 1139 8899 1173
rect 8937 1139 8971 1173
rect 9009 1139 9043 1173
rect 9081 1139 9115 1173
rect 9153 1139 9187 1173
rect 9225 1139 9259 1173
rect 9297 1139 9331 1173
rect 9369 1139 9403 1173
rect 9441 1139 9475 1173
rect 9513 1139 9547 1173
rect 9585 1139 9619 1173
rect 9657 1139 9691 1173
rect 6502 987 6536 1021
rect 6502 915 6536 949
rect 6502 843 6536 877
rect 6502 771 6536 805
rect 6502 699 6536 733
rect 6502 627 6536 661
rect 6502 555 6536 589
rect 6502 483 6536 517
rect 6502 411 6536 445
rect 6502 339 6536 373
rect 6502 267 6536 301
rect 6502 195 6536 229
rect 6502 123 6536 157
rect 6502 51 6536 85
rect 6502 -21 6536 13
rect 6502 -93 6536 -59
rect 6502 -165 6536 -131
rect 6502 -237 6536 -203
rect 6502 -309 6536 -275
rect -92 -1714 -58 -1680
rect -20 -1714 14 -1680
rect 52 -1714 86 -1680
rect 124 -1714 158 -1680
rect 196 -1714 230 -1680
rect 268 -1714 302 -1680
rect 340 -1714 374 -1680
rect 412 -1714 446 -1680
rect 484 -1714 518 -1680
rect 556 -1714 590 -1680
rect 628 -1714 662 -1680
rect 700 -1714 734 -1680
rect 772 -1714 806 -1680
rect 844 -1714 878 -1680
rect 916 -1714 950 -1680
rect 988 -1714 1022 -1680
rect 1060 -1714 1094 -1680
rect 1132 -1714 1166 -1680
rect 1204 -1714 1238 -1680
rect 1276 -1714 1310 -1680
rect 1348 -1714 1382 -1680
rect 1420 -1714 1454 -1680
rect 1492 -1714 1526 -1680
rect 1564 -1714 1598 -1680
rect 1636 -1714 1670 -1680
rect 1708 -1714 1742 -1680
rect 1780 -1714 1814 -1680
rect 1852 -1714 1886 -1680
rect 1924 -1714 1958 -1680
rect 1996 -1714 2030 -1680
rect 2068 -1714 2102 -1680
rect 2140 -1714 2174 -1680
rect 2212 -1714 2246 -1680
rect 2284 -1714 2318 -1680
rect 2356 -1714 2390 -1680
rect 2428 -1714 2462 -1680
rect 2500 -1714 2534 -1680
rect 2572 -1714 2606 -1680
rect 2644 -1714 2678 -1680
rect 2716 -1714 2750 -1680
rect 2788 -1714 2822 -1680
rect 2860 -1714 2894 -1680
rect 2932 -1714 2966 -1680
rect 3004 -1714 3038 -1680
rect 3076 -1714 3110 -1680
rect 3148 -1714 3182 -1680
rect 3220 -1714 3254 -1680
rect 3292 -1714 3326 -1680
rect 3364 -1714 3398 -1680
rect 3436 -1714 3470 -1680
rect 3508 -1714 3542 -1680
rect 3580 -1714 3614 -1680
rect 3652 -1714 3686 -1680
rect 3724 -1714 3758 -1680
rect 3796 -1714 3830 -1680
rect 3868 -1714 3902 -1680
rect 3940 -1714 3974 -1680
rect 4012 -1714 4046 -1680
rect 4084 -1714 4118 -1680
rect 4156 -1714 4190 -1680
rect 4228 -1714 4262 -1680
rect 4300 -1714 4334 -1680
rect 4372 -1714 4406 -1680
rect 4444 -1714 4478 -1680
rect 4516 -1714 4550 -1680
rect 4588 -1714 4622 -1680
rect 4660 -1714 4694 -1680
rect 4732 -1714 4766 -1680
rect 4804 -1714 4838 -1680
rect 4876 -1714 4910 -1680
rect 4948 -1714 4982 -1680
rect 5020 -1714 5054 -1680
rect 5092 -1714 5126 -1680
rect 5164 -1714 5198 -1680
rect 5236 -1714 5270 -1680
rect 5308 -1714 5342 -1680
rect 5380 -1714 5414 -1680
rect 5452 -1714 5486 -1680
rect 5524 -1714 5558 -1680
rect 5596 -1714 5630 -1680
rect 5668 -1714 5702 -1680
rect 5740 -1714 5774 -1680
rect 5812 -1714 5846 -1680
rect 5884 -1714 5918 -1680
rect 5956 -1714 5990 -1680
rect 6028 -1714 6062 -1680
rect 6100 -1714 6134 -1680
rect 6172 -1714 6206 -1680
rect 6244 -1714 6278 -1680
rect 6316 -1714 6350 -1680
rect 6388 -1714 6422 -1680
rect 6460 -1714 6494 -1680
rect 6532 -1714 6566 -1680
rect 6604 -1714 6638 -1680
rect 6676 -1714 6710 -1680
rect 6748 -1714 6782 -1680
rect 6820 -1714 6854 -1680
rect 6892 -1714 6926 -1680
rect 6964 -1714 6998 -1680
rect 7036 -1714 7070 -1680
rect 7108 -1714 7142 -1680
rect 7180 -1714 7214 -1680
rect 7252 -1714 7286 -1680
rect 7324 -1714 7358 -1680
rect 7396 -1714 7430 -1680
rect 7468 -1714 7502 -1680
rect 7540 -1714 7574 -1680
rect 7612 -1714 7646 -1680
rect 7684 -1714 7718 -1680
rect 7756 -1714 7790 -1680
rect 7828 -1714 7862 -1680
rect 7900 -1714 7934 -1680
rect 7972 -1714 8006 -1680
rect 8044 -1714 8078 -1680
rect 8116 -1714 8150 -1680
rect 8188 -1714 8222 -1680
rect 8260 -1714 8294 -1680
rect 8332 -1714 8366 -1680
rect 8404 -1714 8438 -1680
rect 8476 -1714 8510 -1680
rect 8548 -1714 8582 -1680
rect 8620 -1714 8654 -1680
rect 8692 -1714 8726 -1680
rect 8764 -1714 8798 -1680
rect 8836 -1714 8870 -1680
rect 8908 -1714 8942 -1680
rect 8980 -1714 9014 -1680
rect 9052 -1714 9086 -1680
rect 9124 -1714 9158 -1680
rect 9196 -1714 9230 -1680
rect 9268 -1714 9302 -1680
rect 9340 -1714 9374 -1680
rect 9412 -1714 9446 -1680
rect 9484 -1714 9518 -1680
rect 9556 -1714 9590 -1680
rect 9628 -1714 9662 -1680
rect 9700 -1714 9734 -1680
rect 9772 -1714 9806 -1680
rect 9844 -1714 9878 -1680
<< metal1 >>
rect -118 1173 9870 1280
rect -118 1169 61 1173
rect 14 1139 61 1169
rect 95 1139 133 1173
rect 167 1139 205 1173
rect 239 1139 277 1173
rect 311 1139 349 1173
rect 383 1139 421 1173
rect 455 1139 493 1173
rect 527 1139 565 1173
rect 599 1139 637 1173
rect 671 1139 709 1173
rect 743 1139 781 1173
rect 815 1139 853 1173
rect 887 1139 925 1173
rect 959 1139 997 1173
rect 1031 1139 1069 1173
rect 1103 1139 1141 1173
rect 1175 1139 1213 1173
rect 1247 1139 1285 1173
rect 1319 1139 1357 1173
rect 1391 1139 1429 1173
rect 1463 1139 1501 1173
rect 1535 1139 1573 1173
rect 1607 1139 1645 1173
rect 1679 1139 1717 1173
rect 1751 1139 1789 1173
rect 1823 1139 1861 1173
rect 1895 1139 1933 1173
rect 1967 1139 2005 1173
rect 2039 1139 2077 1173
rect 2111 1139 2149 1173
rect 2183 1139 2221 1173
rect 2255 1139 2293 1173
rect 2327 1139 2365 1173
rect 2399 1139 2437 1173
rect 2471 1139 2509 1173
rect 2543 1139 2581 1173
rect 2615 1139 2653 1173
rect 2687 1139 2725 1173
rect 2759 1139 2797 1173
rect 2831 1139 2869 1173
rect 2903 1139 2941 1173
rect 2975 1139 3013 1173
rect 3047 1139 3085 1173
rect 3119 1169 3347 1173
rect 3119 1139 3166 1169
rect 14 1133 3166 1139
rect 3300 1139 3347 1169
rect 3381 1139 3419 1173
rect 3453 1139 3491 1173
rect 3525 1139 3563 1173
rect 3597 1139 3635 1173
rect 3669 1139 3707 1173
rect 3741 1139 3779 1173
rect 3813 1139 3851 1173
rect 3885 1139 3923 1173
rect 3957 1139 3995 1173
rect 4029 1139 4067 1173
rect 4101 1139 4139 1173
rect 4173 1139 4211 1173
rect 4245 1139 4283 1173
rect 4317 1139 4355 1173
rect 4389 1139 4427 1173
rect 4461 1139 4499 1173
rect 4533 1139 4571 1173
rect 4605 1139 4643 1173
rect 4677 1139 4715 1173
rect 4749 1139 4787 1173
rect 4821 1139 4859 1173
rect 4893 1139 4931 1173
rect 4965 1139 5003 1173
rect 5037 1139 5075 1173
rect 5109 1139 5147 1173
rect 5181 1139 5219 1173
rect 5253 1139 5291 1173
rect 5325 1139 5363 1173
rect 5397 1139 5435 1173
rect 5469 1139 5507 1173
rect 5541 1139 5579 1173
rect 5613 1139 5651 1173
rect 5685 1139 5723 1173
rect 5757 1139 5795 1173
rect 5829 1139 5867 1173
rect 5901 1139 5939 1173
rect 5973 1139 6011 1173
rect 6045 1139 6083 1173
rect 6117 1139 6155 1173
rect 6189 1139 6227 1173
rect 6261 1139 6299 1173
rect 6333 1139 6371 1173
rect 6405 1139 6633 1173
rect 6667 1139 6705 1173
rect 6739 1139 6777 1173
rect 6811 1139 6849 1173
rect 6883 1139 6921 1173
rect 6955 1139 6993 1173
rect 7027 1139 7065 1173
rect 7099 1139 7137 1173
rect 7171 1139 7209 1173
rect 7243 1139 7281 1173
rect 7315 1139 7353 1173
rect 7387 1139 7425 1173
rect 7459 1139 7497 1173
rect 7531 1139 7569 1173
rect 7603 1139 7641 1173
rect 7675 1139 7713 1173
rect 7747 1139 7785 1173
rect 7819 1139 7857 1173
rect 7891 1139 7929 1173
rect 7963 1139 8001 1173
rect 8035 1139 8073 1173
rect 8107 1139 8145 1173
rect 8179 1139 8217 1173
rect 8251 1139 8289 1173
rect 8323 1139 8361 1173
rect 8395 1139 8433 1173
rect 8467 1139 8505 1173
rect 8539 1139 8577 1173
rect 8611 1139 8649 1173
rect 8683 1139 8721 1173
rect 8755 1139 8793 1173
rect 8827 1139 8865 1173
rect 8899 1139 8937 1173
rect 8971 1139 9009 1173
rect 9043 1139 9081 1173
rect 9115 1139 9153 1173
rect 9187 1139 9225 1173
rect 9259 1139 9297 1173
rect 9331 1139 9369 1173
rect 9403 1139 9441 1173
rect 9475 1139 9513 1173
rect 9547 1139 9585 1173
rect 9619 1139 9657 1173
rect 9691 1169 9870 1173
rect 9691 1139 9738 1169
rect 3300 1133 9738 1139
rect 3366 1093 6386 1097
rect 3366 1041 3378 1093
rect 3430 1041 3442 1093
rect 3494 1041 3506 1093
rect 3558 1041 3570 1093
rect 3622 1041 3634 1093
rect 3686 1041 3698 1093
rect 3750 1041 3762 1093
rect 3814 1041 3826 1093
rect 3878 1041 3890 1093
rect 3942 1041 3954 1093
rect 4006 1041 4018 1093
rect 4070 1041 4082 1093
rect 4134 1041 4146 1093
rect 4198 1041 4210 1093
rect 4262 1041 4274 1093
rect 4326 1041 4338 1093
rect 4390 1041 4402 1093
rect 4454 1041 4466 1093
rect 4518 1041 4530 1093
rect 4582 1041 4594 1093
rect 4646 1041 4658 1093
rect 4710 1041 4722 1093
rect 4774 1041 4786 1093
rect 4838 1041 4850 1093
rect 4902 1041 4914 1093
rect 4966 1041 4978 1093
rect 5030 1041 5042 1093
rect 5094 1041 5106 1093
rect 5158 1041 5170 1093
rect 5222 1041 5234 1093
rect 5286 1041 5298 1093
rect 5350 1041 5362 1093
rect 5414 1041 5426 1093
rect 5478 1041 5490 1093
rect 5542 1041 5554 1093
rect 5606 1041 5618 1093
rect 5670 1041 5682 1093
rect 5734 1041 5746 1093
rect 5798 1041 5810 1093
rect 5862 1041 5874 1093
rect 5926 1041 5938 1093
rect 5990 1041 6002 1093
rect 6054 1041 6066 1093
rect 6118 1041 6130 1093
rect 6182 1041 6194 1093
rect 6246 1041 6258 1093
rect 6310 1041 6322 1093
rect 6374 1041 6386 1093
rect 3366 1037 6386 1041
rect 6434 1021 6604 1133
rect 6434 987 6502 1021
rect 6536 987 6604 1021
rect 6434 956 6604 987
rect -11 -244 90 956
rect 3080 926 3158 956
rect 3080 874 3093 926
rect 3145 874 3158 926
rect 3080 862 3158 874
rect 3080 810 3093 862
rect 3145 810 3158 862
rect 3080 798 3158 810
rect 3080 746 3093 798
rect 3145 746 3158 798
rect 3080 734 3158 746
rect 3080 682 3093 734
rect 3145 682 3158 734
rect 3080 670 3158 682
rect 3080 618 3093 670
rect 3145 618 3158 670
rect 3080 606 3158 618
rect 3080 554 3093 606
rect 3145 554 3158 606
rect 3080 542 3158 554
rect 3080 490 3093 542
rect 3145 490 3158 542
rect 3080 478 3158 490
rect 3080 426 3093 478
rect 3145 426 3158 478
rect 3080 414 3158 426
rect 3080 362 3093 414
rect 3145 362 3158 414
rect 3080 350 3158 362
rect 3080 298 3093 350
rect 3145 298 3158 350
rect 3080 286 3158 298
rect 3080 234 3093 286
rect 3145 234 3158 286
rect 3080 222 3158 234
rect 3080 170 3093 222
rect 3145 170 3158 222
rect 3080 158 3158 170
rect 3080 106 3093 158
rect 3145 106 3158 158
rect 3080 94 3158 106
rect 3080 42 3093 94
rect 3145 42 3158 94
rect 3080 30 3158 42
rect 3080 -22 3093 30
rect 3145 -22 3158 30
rect 3080 -34 3158 -22
rect 3080 -86 3093 -34
rect 3145 -86 3158 -34
rect 3080 -98 3158 -86
rect 3080 -150 3093 -98
rect 3145 -150 3158 -98
rect 3080 -162 3158 -150
rect 3080 -214 3093 -162
rect 3145 -214 3158 -162
rect 3080 -244 3158 -214
rect 3308 926 3386 956
rect 3308 874 3321 926
rect 3373 874 3386 926
rect 3308 862 3386 874
rect 3308 810 3321 862
rect 3373 810 3386 862
rect 3308 798 3386 810
rect 3308 746 3321 798
rect 3373 746 3386 798
rect 3308 734 3386 746
rect 3308 682 3321 734
rect 3373 682 3386 734
rect 3308 670 3386 682
rect 3308 618 3321 670
rect 3373 618 3386 670
rect 3308 606 3386 618
rect 3308 554 3321 606
rect 3373 554 3386 606
rect 3308 542 3386 554
rect 3308 490 3321 542
rect 3373 490 3386 542
rect 3308 478 3386 490
rect 3308 426 3321 478
rect 3373 426 3386 478
rect 3308 414 3386 426
rect 3308 362 3321 414
rect 3373 362 3386 414
rect 3308 350 3386 362
rect 3308 298 3321 350
rect 3373 298 3386 350
rect 3308 286 3386 298
rect 3308 234 3321 286
rect 3373 234 3386 286
rect 3308 222 3386 234
rect 3308 170 3321 222
rect 3373 170 3386 222
rect 3308 158 3386 170
rect 3308 106 3321 158
rect 3373 106 3386 158
rect 3308 94 3386 106
rect 3308 42 3321 94
rect 3373 42 3386 94
rect 3308 30 3386 42
rect 3308 -22 3321 30
rect 3373 -22 3386 30
rect 3308 -34 3386 -22
rect 3308 -86 3321 -34
rect 3373 -86 3386 -34
rect 3308 -98 3386 -86
rect 3308 -150 3321 -98
rect 3373 -150 3386 -98
rect 3308 -162 3386 -150
rect 3308 -214 3321 -162
rect 3373 -214 3386 -162
rect 3308 -244 3386 -214
rect 6382 949 6656 956
rect 6382 915 6502 949
rect 6536 915 6656 949
rect 6382 877 6656 915
rect 6382 843 6502 877
rect 6536 843 6656 877
rect 6382 805 6656 843
rect 6382 771 6502 805
rect 6536 771 6656 805
rect 6382 733 6656 771
rect 6382 699 6502 733
rect 6536 699 6656 733
rect 6382 661 6656 699
rect 6382 627 6502 661
rect 6536 627 6656 661
rect 6382 589 6656 627
rect 6382 555 6502 589
rect 6536 555 6656 589
rect 6382 517 6656 555
rect 6382 483 6502 517
rect 6536 483 6656 517
rect 6382 445 6656 483
rect 6382 411 6502 445
rect 6536 411 6656 445
rect 6382 373 6656 411
rect 6382 339 6502 373
rect 6536 339 6656 373
rect 6382 301 6656 339
rect 6382 267 6502 301
rect 6536 267 6656 301
rect 6382 229 6656 267
rect 6382 195 6502 229
rect 6536 195 6656 229
rect 6382 157 6656 195
rect 6382 123 6502 157
rect 6536 123 6656 157
rect 6382 85 6656 123
rect 6382 51 6502 85
rect 6536 51 6656 85
rect 6382 13 6656 51
rect 6382 -21 6502 13
rect 6536 -21 6656 13
rect 6382 -59 6656 -21
rect 6382 -93 6502 -59
rect 6536 -93 6656 -59
rect 6382 -131 6656 -93
rect 6382 -165 6502 -131
rect 6536 -165 6656 -131
rect 6382 -203 6656 -165
rect 6382 -237 6502 -203
rect 6536 -237 6656 -203
rect 6382 -244 6656 -237
rect 9662 -244 9761 956
rect -11 -463 39 -244
rect 6496 -275 6542 -244
rect -71 -487 39 -463
rect -71 -539 -37 -487
rect 15 -539 39 -487
rect -71 -563 39 -539
rect -11 -1037 39 -563
rect 93 -727 143 -285
rect 6496 -309 6502 -275
rect 6536 -309 6542 -275
rect 6496 -343 6542 -309
rect 6665 -448 6715 -285
rect 6610 -456 6730 -448
rect 6610 -572 6612 -456
rect 6728 -572 6730 -456
rect 9711 -463 9761 -244
rect 9701 -487 9821 -463
rect 9701 -539 9735 -487
rect 9787 -539 9821 -487
rect 9701 -563 9821 -539
rect 6610 -580 6730 -572
rect 83 -751 203 -727
rect 83 -803 117 -751
rect 169 -803 203 -751
rect 83 -827 203 -803
rect 93 -1005 143 -827
rect 6665 -1005 6715 -580
rect 9711 -1037 9761 -563
rect -11 -1437 89 -1037
rect 3095 -1437 3369 -1037
rect 6365 -1051 6443 -1037
rect 6365 -1103 6378 -1051
rect 6430 -1103 6443 -1051
rect 6365 -1115 6443 -1103
rect 6365 -1167 6378 -1115
rect 6430 -1167 6443 -1115
rect 6365 -1179 6443 -1167
rect 6365 -1231 6378 -1179
rect 6430 -1231 6443 -1179
rect 6365 -1243 6443 -1231
rect 6365 -1295 6378 -1243
rect 6430 -1295 6443 -1243
rect 6365 -1307 6443 -1295
rect 6365 -1359 6378 -1307
rect 6430 -1359 6443 -1307
rect 6365 -1371 6443 -1359
rect 6365 -1423 6378 -1371
rect 6430 -1423 6443 -1371
rect 6365 -1437 6443 -1423
rect 6593 -1051 6671 -1037
rect 6593 -1103 6606 -1051
rect 6658 -1103 6671 -1051
rect 6593 -1115 6671 -1103
rect 6593 -1167 6606 -1115
rect 6658 -1167 6671 -1115
rect 6593 -1179 6671 -1167
rect 6593 -1231 6606 -1179
rect 6658 -1231 6671 -1179
rect 6593 -1243 6671 -1231
rect 6593 -1295 6606 -1243
rect 6658 -1295 6671 -1243
rect 6593 -1307 6671 -1295
rect 6593 -1359 6606 -1307
rect 6658 -1359 6671 -1307
rect 6593 -1371 6671 -1359
rect 6593 -1423 6606 -1371
rect 6658 -1423 6671 -1371
rect 6593 -1437 6671 -1423
rect 9661 -1437 9761 -1037
rect 3147 -1641 3317 -1437
rect 3365 -1513 6385 -1509
rect 3365 -1565 3377 -1513
rect 3429 -1565 3441 -1513
rect 3493 -1565 3505 -1513
rect 3557 -1565 3569 -1513
rect 3621 -1565 3633 -1513
rect 3685 -1565 3697 -1513
rect 3749 -1565 3761 -1513
rect 3813 -1565 3825 -1513
rect 3877 -1565 3889 -1513
rect 3941 -1565 3953 -1513
rect 4005 -1565 4017 -1513
rect 4069 -1565 4081 -1513
rect 4133 -1565 4145 -1513
rect 4197 -1565 4209 -1513
rect 4261 -1565 4273 -1513
rect 4325 -1565 4337 -1513
rect 4389 -1565 4401 -1513
rect 4453 -1565 4465 -1513
rect 4517 -1565 4529 -1513
rect 4581 -1565 4593 -1513
rect 4645 -1565 4657 -1513
rect 4709 -1565 4721 -1513
rect 4773 -1565 4785 -1513
rect 4837 -1565 4849 -1513
rect 4901 -1565 4913 -1513
rect 4965 -1565 4977 -1513
rect 5029 -1565 5041 -1513
rect 5093 -1565 5105 -1513
rect 5157 -1565 5169 -1513
rect 5221 -1565 5233 -1513
rect 5285 -1565 5297 -1513
rect 5349 -1565 5361 -1513
rect 5413 -1565 5425 -1513
rect 5477 -1565 5489 -1513
rect 5541 -1565 5553 -1513
rect 5605 -1565 5617 -1513
rect 5669 -1565 5681 -1513
rect 5733 -1565 5745 -1513
rect 5797 -1565 5809 -1513
rect 5861 -1565 5873 -1513
rect 5925 -1565 5937 -1513
rect 5989 -1565 6001 -1513
rect 6053 -1565 6065 -1513
rect 6117 -1565 6129 -1513
rect 6181 -1565 6193 -1513
rect 6245 -1565 6257 -1513
rect 6309 -1565 6321 -1513
rect 6373 -1565 6385 -1513
rect 3365 -1569 6385 -1565
rect -119 -1680 9905 -1641
rect -119 -1714 -92 -1680
rect -58 -1714 -20 -1680
rect 14 -1714 52 -1680
rect 86 -1714 124 -1680
rect 158 -1714 196 -1680
rect 230 -1714 268 -1680
rect 302 -1714 340 -1680
rect 374 -1714 412 -1680
rect 446 -1714 484 -1680
rect 518 -1714 556 -1680
rect 590 -1714 628 -1680
rect 662 -1714 700 -1680
rect 734 -1714 772 -1680
rect 806 -1714 844 -1680
rect 878 -1714 916 -1680
rect 950 -1714 988 -1680
rect 1022 -1714 1060 -1680
rect 1094 -1714 1132 -1680
rect 1166 -1714 1204 -1680
rect 1238 -1714 1276 -1680
rect 1310 -1714 1348 -1680
rect 1382 -1714 1420 -1680
rect 1454 -1714 1492 -1680
rect 1526 -1714 1564 -1680
rect 1598 -1714 1636 -1680
rect 1670 -1714 1708 -1680
rect 1742 -1714 1780 -1680
rect 1814 -1714 1852 -1680
rect 1886 -1714 1924 -1680
rect 1958 -1714 1996 -1680
rect 2030 -1714 2068 -1680
rect 2102 -1714 2140 -1680
rect 2174 -1714 2212 -1680
rect 2246 -1714 2284 -1680
rect 2318 -1714 2356 -1680
rect 2390 -1714 2428 -1680
rect 2462 -1714 2500 -1680
rect 2534 -1714 2572 -1680
rect 2606 -1714 2644 -1680
rect 2678 -1714 2716 -1680
rect 2750 -1714 2788 -1680
rect 2822 -1714 2860 -1680
rect 2894 -1714 2932 -1680
rect 2966 -1714 3004 -1680
rect 3038 -1714 3076 -1680
rect 3110 -1714 3148 -1680
rect 3182 -1714 3220 -1680
rect 3254 -1714 3292 -1680
rect 3326 -1714 3364 -1680
rect 3398 -1714 3436 -1680
rect 3470 -1714 3508 -1680
rect 3542 -1714 3580 -1680
rect 3614 -1714 3652 -1680
rect 3686 -1714 3724 -1680
rect 3758 -1714 3796 -1680
rect 3830 -1714 3868 -1680
rect 3902 -1714 3940 -1680
rect 3974 -1714 4012 -1680
rect 4046 -1714 4084 -1680
rect 4118 -1714 4156 -1680
rect 4190 -1714 4228 -1680
rect 4262 -1714 4300 -1680
rect 4334 -1714 4372 -1680
rect 4406 -1714 4444 -1680
rect 4478 -1714 4516 -1680
rect 4550 -1714 4588 -1680
rect 4622 -1714 4660 -1680
rect 4694 -1714 4732 -1680
rect 4766 -1714 4804 -1680
rect 4838 -1714 4876 -1680
rect 4910 -1714 4948 -1680
rect 4982 -1714 5020 -1680
rect 5054 -1714 5092 -1680
rect 5126 -1714 5164 -1680
rect 5198 -1714 5236 -1680
rect 5270 -1714 5308 -1680
rect 5342 -1714 5380 -1680
rect 5414 -1714 5452 -1680
rect 5486 -1714 5524 -1680
rect 5558 -1714 5596 -1680
rect 5630 -1714 5668 -1680
rect 5702 -1714 5740 -1680
rect 5774 -1714 5812 -1680
rect 5846 -1714 5884 -1680
rect 5918 -1714 5956 -1680
rect 5990 -1714 6028 -1680
rect 6062 -1714 6100 -1680
rect 6134 -1714 6172 -1680
rect 6206 -1714 6244 -1680
rect 6278 -1714 6316 -1680
rect 6350 -1714 6388 -1680
rect 6422 -1714 6460 -1680
rect 6494 -1714 6532 -1680
rect 6566 -1714 6604 -1680
rect 6638 -1714 6676 -1680
rect 6710 -1714 6748 -1680
rect 6782 -1714 6820 -1680
rect 6854 -1714 6892 -1680
rect 6926 -1714 6964 -1680
rect 6998 -1714 7036 -1680
rect 7070 -1714 7108 -1680
rect 7142 -1714 7180 -1680
rect 7214 -1714 7252 -1680
rect 7286 -1714 7324 -1680
rect 7358 -1714 7396 -1680
rect 7430 -1714 7468 -1680
rect 7502 -1714 7540 -1680
rect 7574 -1714 7612 -1680
rect 7646 -1714 7684 -1680
rect 7718 -1714 7756 -1680
rect 7790 -1714 7828 -1680
rect 7862 -1714 7900 -1680
rect 7934 -1714 7972 -1680
rect 8006 -1714 8044 -1680
rect 8078 -1714 8116 -1680
rect 8150 -1714 8188 -1680
rect 8222 -1714 8260 -1680
rect 8294 -1714 8332 -1680
rect 8366 -1714 8404 -1680
rect 8438 -1714 8476 -1680
rect 8510 -1714 8548 -1680
rect 8582 -1714 8620 -1680
rect 8654 -1714 8692 -1680
rect 8726 -1714 8764 -1680
rect 8798 -1714 8836 -1680
rect 8870 -1714 8908 -1680
rect 8942 -1714 8980 -1680
rect 9014 -1714 9052 -1680
rect 9086 -1714 9124 -1680
rect 9158 -1714 9196 -1680
rect 9230 -1714 9268 -1680
rect 9302 -1714 9340 -1680
rect 9374 -1714 9412 -1680
rect 9446 -1714 9484 -1680
rect 9518 -1714 9556 -1680
rect 9590 -1714 9628 -1680
rect 9662 -1714 9700 -1680
rect 9734 -1714 9772 -1680
rect 9806 -1714 9844 -1680
rect 9878 -1714 9905 -1680
rect -119 -1753 9905 -1714
<< via1 >>
rect 3378 1041 3430 1093
rect 3442 1041 3494 1093
rect 3506 1041 3558 1093
rect 3570 1041 3622 1093
rect 3634 1041 3686 1093
rect 3698 1041 3750 1093
rect 3762 1041 3814 1093
rect 3826 1041 3878 1093
rect 3890 1041 3942 1093
rect 3954 1041 4006 1093
rect 4018 1041 4070 1093
rect 4082 1041 4134 1093
rect 4146 1041 4198 1093
rect 4210 1041 4262 1093
rect 4274 1041 4326 1093
rect 4338 1041 4390 1093
rect 4402 1041 4454 1093
rect 4466 1041 4518 1093
rect 4530 1041 4582 1093
rect 4594 1041 4646 1093
rect 4658 1041 4710 1093
rect 4722 1041 4774 1093
rect 4786 1041 4838 1093
rect 4850 1041 4902 1093
rect 4914 1041 4966 1093
rect 4978 1041 5030 1093
rect 5042 1041 5094 1093
rect 5106 1041 5158 1093
rect 5170 1041 5222 1093
rect 5234 1041 5286 1093
rect 5298 1041 5350 1093
rect 5362 1041 5414 1093
rect 5426 1041 5478 1093
rect 5490 1041 5542 1093
rect 5554 1041 5606 1093
rect 5618 1041 5670 1093
rect 5682 1041 5734 1093
rect 5746 1041 5798 1093
rect 5810 1041 5862 1093
rect 5874 1041 5926 1093
rect 5938 1041 5990 1093
rect 6002 1041 6054 1093
rect 6066 1041 6118 1093
rect 6130 1041 6182 1093
rect 6194 1041 6246 1093
rect 6258 1041 6310 1093
rect 6322 1041 6374 1093
rect 3093 874 3145 926
rect 3093 810 3145 862
rect 3093 746 3145 798
rect 3093 682 3145 734
rect 3093 618 3145 670
rect 3093 554 3145 606
rect 3093 490 3145 542
rect 3093 426 3145 478
rect 3093 362 3145 414
rect 3093 298 3145 350
rect 3093 234 3145 286
rect 3093 170 3145 222
rect 3093 106 3145 158
rect 3093 42 3145 94
rect 3093 -22 3145 30
rect 3093 -86 3145 -34
rect 3093 -150 3145 -98
rect 3093 -214 3145 -162
rect 3321 874 3373 926
rect 3321 810 3373 862
rect 3321 746 3373 798
rect 3321 682 3373 734
rect 3321 618 3373 670
rect 3321 554 3373 606
rect 3321 490 3373 542
rect 3321 426 3373 478
rect 3321 362 3373 414
rect 3321 298 3373 350
rect 3321 234 3373 286
rect 3321 170 3373 222
rect 3321 106 3373 158
rect 3321 42 3373 94
rect 3321 -22 3373 30
rect 3321 -86 3373 -34
rect 3321 -150 3373 -98
rect 3321 -214 3373 -162
rect -37 -539 15 -487
rect 6612 -572 6728 -456
rect 9735 -539 9787 -487
rect 117 -803 169 -751
rect 6378 -1103 6430 -1051
rect 6378 -1167 6430 -1115
rect 6378 -1231 6430 -1179
rect 6378 -1295 6430 -1243
rect 6378 -1359 6430 -1307
rect 6378 -1423 6430 -1371
rect 6606 -1103 6658 -1051
rect 6606 -1167 6658 -1115
rect 6606 -1231 6658 -1179
rect 6606 -1295 6658 -1243
rect 6606 -1359 6658 -1307
rect 6606 -1423 6658 -1371
rect 3377 -1565 3429 -1513
rect 3441 -1565 3493 -1513
rect 3505 -1565 3557 -1513
rect 3569 -1565 3621 -1513
rect 3633 -1565 3685 -1513
rect 3697 -1565 3749 -1513
rect 3761 -1565 3813 -1513
rect 3825 -1565 3877 -1513
rect 3889 -1565 3941 -1513
rect 3953 -1565 4005 -1513
rect 4017 -1565 4069 -1513
rect 4081 -1565 4133 -1513
rect 4145 -1565 4197 -1513
rect 4209 -1565 4261 -1513
rect 4273 -1565 4325 -1513
rect 4337 -1565 4389 -1513
rect 4401 -1565 4453 -1513
rect 4465 -1565 4517 -1513
rect 4529 -1565 4581 -1513
rect 4593 -1565 4645 -1513
rect 4657 -1565 4709 -1513
rect 4721 -1565 4773 -1513
rect 4785 -1565 4837 -1513
rect 4849 -1565 4901 -1513
rect 4913 -1565 4965 -1513
rect 4977 -1565 5029 -1513
rect 5041 -1565 5093 -1513
rect 5105 -1565 5157 -1513
rect 5169 -1565 5221 -1513
rect 5233 -1565 5285 -1513
rect 5297 -1565 5349 -1513
rect 5361 -1565 5413 -1513
rect 5425 -1565 5477 -1513
rect 5489 -1565 5541 -1513
rect 5553 -1565 5605 -1513
rect 5617 -1565 5669 -1513
rect 5681 -1565 5733 -1513
rect 5745 -1565 5797 -1513
rect 5809 -1565 5861 -1513
rect 5873 -1565 5925 -1513
rect 5937 -1565 5989 -1513
rect 6001 -1565 6053 -1513
rect 6065 -1565 6117 -1513
rect 6129 -1565 6181 -1513
rect 6193 -1565 6245 -1513
rect 6257 -1565 6309 -1513
rect 6321 -1565 6373 -1513
<< metal2 >>
rect -106 1093 6376 1107
rect -106 1041 3378 1093
rect 3430 1041 3442 1093
rect 3494 1041 3506 1093
rect 3558 1041 3570 1093
rect 3622 1041 3634 1093
rect 3686 1041 3698 1093
rect 3750 1041 3762 1093
rect 3814 1041 3826 1093
rect 3878 1041 3890 1093
rect 3942 1041 3954 1093
rect 4006 1041 4018 1093
rect 4070 1041 4082 1093
rect 4134 1041 4146 1093
rect 4198 1041 4210 1093
rect 4262 1041 4274 1093
rect 4326 1041 4338 1093
rect 4390 1041 4402 1093
rect 4454 1041 4466 1093
rect 4518 1041 4530 1093
rect 4582 1041 4594 1093
rect 4646 1041 4658 1093
rect 4710 1041 4722 1093
rect 4774 1041 4786 1093
rect 4838 1041 4850 1093
rect 4902 1041 4914 1093
rect 4966 1041 4978 1093
rect 5030 1041 5042 1093
rect 5094 1041 5106 1093
rect 5158 1041 5170 1093
rect 5222 1041 5234 1093
rect 5286 1041 5298 1093
rect 5350 1041 5362 1093
rect 5414 1041 5426 1093
rect 5478 1041 5490 1093
rect 5542 1041 5554 1093
rect 5606 1041 5618 1093
rect 5670 1041 5682 1093
rect 5734 1041 5746 1093
rect 5798 1041 5810 1093
rect 5862 1041 5874 1093
rect 5926 1041 5938 1093
rect 5990 1041 6002 1093
rect 6054 1041 6066 1093
rect 6118 1041 6130 1093
rect 6182 1041 6194 1093
rect 6246 1041 6258 1093
rect 6310 1041 6322 1093
rect 6374 1041 6376 1093
rect -106 1027 6376 1041
rect 3090 926 3376 966
rect 3090 874 3093 926
rect 3145 874 3321 926
rect 3373 874 3376 926
rect 3090 862 3376 874
rect 3090 810 3093 862
rect 3145 810 3321 862
rect 3373 810 3376 862
rect 3090 798 3376 810
rect 3090 746 3093 798
rect 3145 746 3321 798
rect 3373 746 3376 798
rect 3090 734 3376 746
rect 3090 682 3093 734
rect 3145 682 3321 734
rect 3373 682 3376 734
rect 3090 670 3376 682
rect 3090 618 3093 670
rect 3145 618 3321 670
rect 3373 618 3376 670
rect 3090 606 3376 618
rect 3090 554 3093 606
rect 3145 554 3321 606
rect 3373 554 3376 606
rect 3090 542 3376 554
rect 3090 490 3093 542
rect 3145 490 3321 542
rect 3373 490 3376 542
rect 3090 478 3376 490
rect 3090 426 3093 478
rect 3145 426 3321 478
rect 3373 426 3376 478
rect 3090 414 3376 426
rect 3090 362 3093 414
rect 3145 362 3321 414
rect 3373 362 3376 414
rect 3090 350 3376 362
rect 3090 298 3093 350
rect 3145 298 3321 350
rect 3373 298 3376 350
rect 3090 286 3376 298
rect 3090 234 3093 286
rect 3145 234 3321 286
rect 3373 234 3376 286
rect 3090 222 3376 234
rect 3090 170 3093 222
rect 3145 170 3321 222
rect 3373 170 3376 222
rect 3090 158 3376 170
rect 3090 106 3093 158
rect 3145 106 3321 158
rect 3373 106 3376 158
rect 3090 94 3376 106
rect 3090 42 3093 94
rect 3145 42 3321 94
rect 3373 42 3376 94
rect 3090 30 3376 42
rect 3090 -22 3093 30
rect 3145 -22 3321 30
rect 3373 -22 3376 30
rect 3090 -34 3376 -22
rect 3090 -86 3093 -34
rect 3145 -86 3321 -34
rect 3373 -86 3376 -34
rect 3090 -98 3376 -86
rect 3090 -150 3093 -98
rect 3145 -150 3321 -98
rect 3373 -150 3376 -98
rect 3090 -162 3376 -150
rect 3090 -214 3093 -162
rect 3145 -214 3321 -162
rect 3373 -214 3376 -162
rect 3090 -254 3376 -214
rect -61 -454 39 -453
rect 6616 -454 6715 -453
rect -62 -456 6736 -454
rect -62 -487 6612 -456
rect -62 -539 -37 -487
rect 15 -539 6612 -487
rect -62 -572 6612 -539
rect 6728 -572 6736 -456
rect -62 -574 6736 -572
rect 9711 -487 9858 -453
rect 9711 -539 9735 -487
rect 9787 -539 9858 -487
rect 9711 -573 9858 -539
rect -107 -751 193 -717
rect -107 -803 117 -751
rect 169 -803 193 -751
rect -107 -837 193 -803
rect 6375 -1051 6661 -1027
rect 6375 -1103 6378 -1051
rect 6430 -1103 6606 -1051
rect 6658 -1103 6661 -1051
rect 6375 -1115 6661 -1103
rect 6375 -1167 6378 -1115
rect 6430 -1167 6606 -1115
rect 6658 -1167 6661 -1115
rect 6375 -1179 6661 -1167
rect 6375 -1231 6378 -1179
rect 6430 -1231 6606 -1179
rect 6658 -1231 6661 -1179
rect 6375 -1243 6661 -1231
rect 6375 -1295 6378 -1243
rect 6430 -1295 6606 -1243
rect 6658 -1295 6661 -1243
rect 6375 -1307 6661 -1295
rect 6375 -1359 6378 -1307
rect 6430 -1359 6606 -1307
rect 6658 -1359 6661 -1307
rect 6375 -1371 6661 -1359
rect 6375 -1423 6378 -1371
rect 6430 -1423 6606 -1371
rect 6658 -1423 6661 -1371
rect 6375 -1447 6661 -1423
rect -107 -1513 6375 -1499
rect -107 -1565 3377 -1513
rect 3429 -1565 3441 -1513
rect 3493 -1565 3505 -1513
rect 3557 -1565 3569 -1513
rect 3621 -1565 3633 -1513
rect 3685 -1565 3697 -1513
rect 3749 -1565 3761 -1513
rect 3813 -1565 3825 -1513
rect 3877 -1565 3889 -1513
rect 3941 -1565 3953 -1513
rect 4005 -1565 4017 -1513
rect 4069 -1565 4081 -1513
rect 4133 -1565 4145 -1513
rect 4197 -1565 4209 -1513
rect 4261 -1565 4273 -1513
rect 4325 -1565 4337 -1513
rect 4389 -1565 4401 -1513
rect 4453 -1565 4465 -1513
rect 4517 -1565 4529 -1513
rect 4581 -1565 4593 -1513
rect 4645 -1565 4657 -1513
rect 4709 -1565 4721 -1513
rect 4773 -1565 4785 -1513
rect 4837 -1565 4849 -1513
rect 4901 -1565 4913 -1513
rect 4965 -1565 4977 -1513
rect 5029 -1565 5041 -1513
rect 5093 -1565 5105 -1513
rect 5157 -1565 5169 -1513
rect 5221 -1565 5233 -1513
rect 5285 -1565 5297 -1513
rect 5349 -1565 5361 -1513
rect 5413 -1565 5425 -1513
rect 5477 -1565 5489 -1513
rect 5541 -1565 5553 -1513
rect 5605 -1565 5617 -1513
rect 5669 -1565 5681 -1513
rect 5733 -1565 5745 -1513
rect 5797 -1565 5809 -1513
rect 5861 -1565 5873 -1513
rect 5925 -1565 5937 -1513
rect 5989 -1565 6001 -1513
rect 6053 -1565 6065 -1513
rect 6117 -1565 6129 -1513
rect 6181 -1565 6193 -1513
rect 6245 -1565 6257 -1513
rect 6309 -1565 6321 -1513
rect 6373 -1565 6375 -1513
rect -107 -1579 6375 -1565
use sky130_fd_pr__pfet_01v8_lvt_NZTZAV  XM1
timestamp 1731265361
transform 1 0 1590 0 1 356
box -1696 -819 1696 819
use sky130_fd_pr__pfet_01v8_lvt_NZTZAV  XM2
timestamp 1731265361
transform 1 0 4876 0 1 356
box -1696 -819 1696 819
use sky130_fd_pr__nfet_01v8_lvt_PHPD3W  XM3
timestamp 1731265361
transform 1 0 1589 0 1 -1237
box -1686 -400 1686 400
use sky130_fd_pr__pfet_01v8_lvt_NZTZAV  XM6
timestamp 1731265361
transform 1 0 8162 0 1 356
box -1696 -819 1696 819
use sky130_fd_pr__nfet_01v8_lvt_PHPD3W  XM7
timestamp 1731265361
transform 1 0 4875 0 1 -1237
box -1686 -400 1686 400
use sky130_fd_pr__nfet_01v8_lvt_PHPD3W  XM8
timestamp 1731265361
transform 1 0 8161 0 1 -1237
box -1686 -400 1686 400
<< labels >>
flabel metal1 s -118 1169 -7 1280 0 FreeSans 1000 0 0 0 VDD
port 1 nsew
flabel metal1 s -107 -1747 -7 -1647 0 FreeSans 1000 0 0 0 VSS
port 2 nsew
flabel metal2 s -42 1027 38 1107 0 FreeSans 1000 0 0 0 VIP
port 3 nsew
flabel metal2 s -38 -1579 42 -1499 0 FreeSans 1000 0 0 0 VIN
port 4 nsew
flabel metal1 s 9711 -687 9761 -637 0 FreeSans 1000 0 0 0 OUT
port 5 nsew
flabel metal2 s -107 -837 13 -717 0 FreeSans 1000 0 0 0 IN
port 6 nsew
<< end >>
