magic
tech sky130A
magscale 1 2
timestamp 1730269323
<< metal3 >>
rect -386 45932 386 45960
rect -386 45508 302 45932
rect 366 45508 386 45932
rect -386 45480 386 45508
rect -386 45212 386 45240
rect -386 44788 302 45212
rect 366 44788 386 45212
rect -386 44760 386 44788
rect -386 44492 386 44520
rect -386 44068 302 44492
rect 366 44068 386 44492
rect -386 44040 386 44068
rect -386 43772 386 43800
rect -386 43348 302 43772
rect 366 43348 386 43772
rect -386 43320 386 43348
rect -386 43052 386 43080
rect -386 42628 302 43052
rect 366 42628 386 43052
rect -386 42600 386 42628
rect -386 42332 386 42360
rect -386 41908 302 42332
rect 366 41908 386 42332
rect -386 41880 386 41908
rect -386 41612 386 41640
rect -386 41188 302 41612
rect 366 41188 386 41612
rect -386 41160 386 41188
rect -386 40892 386 40920
rect -386 40468 302 40892
rect 366 40468 386 40892
rect -386 40440 386 40468
rect -386 40172 386 40200
rect -386 39748 302 40172
rect 366 39748 386 40172
rect -386 39720 386 39748
rect -386 39452 386 39480
rect -386 39028 302 39452
rect 366 39028 386 39452
rect -386 39000 386 39028
rect -386 38732 386 38760
rect -386 38308 302 38732
rect 366 38308 386 38732
rect -386 38280 386 38308
rect -386 38012 386 38040
rect -386 37588 302 38012
rect 366 37588 386 38012
rect -386 37560 386 37588
rect -386 37292 386 37320
rect -386 36868 302 37292
rect 366 36868 386 37292
rect -386 36840 386 36868
rect -386 36572 386 36600
rect -386 36148 302 36572
rect 366 36148 386 36572
rect -386 36120 386 36148
rect -386 35852 386 35880
rect -386 35428 302 35852
rect 366 35428 386 35852
rect -386 35400 386 35428
rect -386 35132 386 35160
rect -386 34708 302 35132
rect 366 34708 386 35132
rect -386 34680 386 34708
rect -386 34412 386 34440
rect -386 33988 302 34412
rect 366 33988 386 34412
rect -386 33960 386 33988
rect -386 33692 386 33720
rect -386 33268 302 33692
rect 366 33268 386 33692
rect -386 33240 386 33268
rect -386 32972 386 33000
rect -386 32548 302 32972
rect 366 32548 386 32972
rect -386 32520 386 32548
rect -386 32252 386 32280
rect -386 31828 302 32252
rect 366 31828 386 32252
rect -386 31800 386 31828
rect -386 31532 386 31560
rect -386 31108 302 31532
rect 366 31108 386 31532
rect -386 31080 386 31108
rect -386 30812 386 30840
rect -386 30388 302 30812
rect 366 30388 386 30812
rect -386 30360 386 30388
rect -386 30092 386 30120
rect -386 29668 302 30092
rect 366 29668 386 30092
rect -386 29640 386 29668
rect -386 29372 386 29400
rect -386 28948 302 29372
rect 366 28948 386 29372
rect -386 28920 386 28948
rect -386 28652 386 28680
rect -386 28228 302 28652
rect 366 28228 386 28652
rect -386 28200 386 28228
rect -386 27932 386 27960
rect -386 27508 302 27932
rect 366 27508 386 27932
rect -386 27480 386 27508
rect -386 27212 386 27240
rect -386 26788 302 27212
rect 366 26788 386 27212
rect -386 26760 386 26788
rect -386 26492 386 26520
rect -386 26068 302 26492
rect 366 26068 386 26492
rect -386 26040 386 26068
rect -386 25772 386 25800
rect -386 25348 302 25772
rect 366 25348 386 25772
rect -386 25320 386 25348
rect -386 25052 386 25080
rect -386 24628 302 25052
rect 366 24628 386 25052
rect -386 24600 386 24628
rect -386 24332 386 24360
rect -386 23908 302 24332
rect 366 23908 386 24332
rect -386 23880 386 23908
rect -386 23612 386 23640
rect -386 23188 302 23612
rect 366 23188 386 23612
rect -386 23160 386 23188
rect -386 22892 386 22920
rect -386 22468 302 22892
rect 366 22468 386 22892
rect -386 22440 386 22468
rect -386 22172 386 22200
rect -386 21748 302 22172
rect 366 21748 386 22172
rect -386 21720 386 21748
rect -386 21452 386 21480
rect -386 21028 302 21452
rect 366 21028 386 21452
rect -386 21000 386 21028
rect -386 20732 386 20760
rect -386 20308 302 20732
rect 366 20308 386 20732
rect -386 20280 386 20308
rect -386 20012 386 20040
rect -386 19588 302 20012
rect 366 19588 386 20012
rect -386 19560 386 19588
rect -386 19292 386 19320
rect -386 18868 302 19292
rect 366 18868 386 19292
rect -386 18840 386 18868
rect -386 18572 386 18600
rect -386 18148 302 18572
rect 366 18148 386 18572
rect -386 18120 386 18148
rect -386 17852 386 17880
rect -386 17428 302 17852
rect 366 17428 386 17852
rect -386 17400 386 17428
rect -386 17132 386 17160
rect -386 16708 302 17132
rect 366 16708 386 17132
rect -386 16680 386 16708
rect -386 16412 386 16440
rect -386 15988 302 16412
rect 366 15988 386 16412
rect -386 15960 386 15988
rect -386 15692 386 15720
rect -386 15268 302 15692
rect 366 15268 386 15692
rect -386 15240 386 15268
rect -386 14972 386 15000
rect -386 14548 302 14972
rect 366 14548 386 14972
rect -386 14520 386 14548
rect -386 14252 386 14280
rect -386 13828 302 14252
rect 366 13828 386 14252
rect -386 13800 386 13828
rect -386 13532 386 13560
rect -386 13108 302 13532
rect 366 13108 386 13532
rect -386 13080 386 13108
rect -386 12812 386 12840
rect -386 12388 302 12812
rect 366 12388 386 12812
rect -386 12360 386 12388
rect -386 12092 386 12120
rect -386 11668 302 12092
rect 366 11668 386 12092
rect -386 11640 386 11668
rect -386 11372 386 11400
rect -386 10948 302 11372
rect 366 10948 386 11372
rect -386 10920 386 10948
rect -386 10652 386 10680
rect -386 10228 302 10652
rect 366 10228 386 10652
rect -386 10200 386 10228
rect -386 9932 386 9960
rect -386 9508 302 9932
rect 366 9508 386 9932
rect -386 9480 386 9508
rect -386 9212 386 9240
rect -386 8788 302 9212
rect 366 8788 386 9212
rect -386 8760 386 8788
rect -386 8492 386 8520
rect -386 8068 302 8492
rect 366 8068 386 8492
rect -386 8040 386 8068
rect -386 7772 386 7800
rect -386 7348 302 7772
rect 366 7348 386 7772
rect -386 7320 386 7348
rect -386 7052 386 7080
rect -386 6628 302 7052
rect 366 6628 386 7052
rect -386 6600 386 6628
rect -386 6332 386 6360
rect -386 5908 302 6332
rect 366 5908 386 6332
rect -386 5880 386 5908
rect -386 5612 386 5640
rect -386 5188 302 5612
rect 366 5188 386 5612
rect -386 5160 386 5188
rect -386 4892 386 4920
rect -386 4468 302 4892
rect 366 4468 386 4892
rect -386 4440 386 4468
rect -386 4172 386 4200
rect -386 3748 302 4172
rect 366 3748 386 4172
rect -386 3720 386 3748
rect -386 3452 386 3480
rect -386 3028 302 3452
rect 366 3028 386 3452
rect -386 3000 386 3028
rect -386 2732 386 2760
rect -386 2308 302 2732
rect 366 2308 386 2732
rect -386 2280 386 2308
rect -386 2012 386 2040
rect -386 1588 302 2012
rect 366 1588 386 2012
rect -386 1560 386 1588
rect -386 1292 386 1320
rect -386 868 302 1292
rect 366 868 386 1292
rect -386 840 386 868
rect -386 572 386 600
rect -386 148 302 572
rect 366 148 386 572
rect -386 120 386 148
rect -386 -148 386 -120
rect -386 -572 302 -148
rect 366 -572 386 -148
rect -386 -600 386 -572
rect -386 -868 386 -840
rect -386 -1292 302 -868
rect 366 -1292 386 -868
rect -386 -1320 386 -1292
rect -386 -1588 386 -1560
rect -386 -2012 302 -1588
rect 366 -2012 386 -1588
rect -386 -2040 386 -2012
rect -386 -2308 386 -2280
rect -386 -2732 302 -2308
rect 366 -2732 386 -2308
rect -386 -2760 386 -2732
rect -386 -3028 386 -3000
rect -386 -3452 302 -3028
rect 366 -3452 386 -3028
rect -386 -3480 386 -3452
rect -386 -3748 386 -3720
rect -386 -4172 302 -3748
rect 366 -4172 386 -3748
rect -386 -4200 386 -4172
rect -386 -4468 386 -4440
rect -386 -4892 302 -4468
rect 366 -4892 386 -4468
rect -386 -4920 386 -4892
rect -386 -5188 386 -5160
rect -386 -5612 302 -5188
rect 366 -5612 386 -5188
rect -386 -5640 386 -5612
rect -386 -5908 386 -5880
rect -386 -6332 302 -5908
rect 366 -6332 386 -5908
rect -386 -6360 386 -6332
rect -386 -6628 386 -6600
rect -386 -7052 302 -6628
rect 366 -7052 386 -6628
rect -386 -7080 386 -7052
rect -386 -7348 386 -7320
rect -386 -7772 302 -7348
rect 366 -7772 386 -7348
rect -386 -7800 386 -7772
rect -386 -8068 386 -8040
rect -386 -8492 302 -8068
rect 366 -8492 386 -8068
rect -386 -8520 386 -8492
rect -386 -8788 386 -8760
rect -386 -9212 302 -8788
rect 366 -9212 386 -8788
rect -386 -9240 386 -9212
rect -386 -9508 386 -9480
rect -386 -9932 302 -9508
rect 366 -9932 386 -9508
rect -386 -9960 386 -9932
rect -386 -10228 386 -10200
rect -386 -10652 302 -10228
rect 366 -10652 386 -10228
rect -386 -10680 386 -10652
rect -386 -10948 386 -10920
rect -386 -11372 302 -10948
rect 366 -11372 386 -10948
rect -386 -11400 386 -11372
rect -386 -11668 386 -11640
rect -386 -12092 302 -11668
rect 366 -12092 386 -11668
rect -386 -12120 386 -12092
rect -386 -12388 386 -12360
rect -386 -12812 302 -12388
rect 366 -12812 386 -12388
rect -386 -12840 386 -12812
rect -386 -13108 386 -13080
rect -386 -13532 302 -13108
rect 366 -13532 386 -13108
rect -386 -13560 386 -13532
rect -386 -13828 386 -13800
rect -386 -14252 302 -13828
rect 366 -14252 386 -13828
rect -386 -14280 386 -14252
rect -386 -14548 386 -14520
rect -386 -14972 302 -14548
rect 366 -14972 386 -14548
rect -386 -15000 386 -14972
rect -386 -15268 386 -15240
rect -386 -15692 302 -15268
rect 366 -15692 386 -15268
rect -386 -15720 386 -15692
rect -386 -15988 386 -15960
rect -386 -16412 302 -15988
rect 366 -16412 386 -15988
rect -386 -16440 386 -16412
rect -386 -16708 386 -16680
rect -386 -17132 302 -16708
rect 366 -17132 386 -16708
rect -386 -17160 386 -17132
rect -386 -17428 386 -17400
rect -386 -17852 302 -17428
rect 366 -17852 386 -17428
rect -386 -17880 386 -17852
rect -386 -18148 386 -18120
rect -386 -18572 302 -18148
rect 366 -18572 386 -18148
rect -386 -18600 386 -18572
rect -386 -18868 386 -18840
rect -386 -19292 302 -18868
rect 366 -19292 386 -18868
rect -386 -19320 386 -19292
rect -386 -19588 386 -19560
rect -386 -20012 302 -19588
rect 366 -20012 386 -19588
rect -386 -20040 386 -20012
rect -386 -20308 386 -20280
rect -386 -20732 302 -20308
rect 366 -20732 386 -20308
rect -386 -20760 386 -20732
rect -386 -21028 386 -21000
rect -386 -21452 302 -21028
rect 366 -21452 386 -21028
rect -386 -21480 386 -21452
rect -386 -21748 386 -21720
rect -386 -22172 302 -21748
rect 366 -22172 386 -21748
rect -386 -22200 386 -22172
rect -386 -22468 386 -22440
rect -386 -22892 302 -22468
rect 366 -22892 386 -22468
rect -386 -22920 386 -22892
rect -386 -23188 386 -23160
rect -386 -23612 302 -23188
rect 366 -23612 386 -23188
rect -386 -23640 386 -23612
rect -386 -23908 386 -23880
rect -386 -24332 302 -23908
rect 366 -24332 386 -23908
rect -386 -24360 386 -24332
rect -386 -24628 386 -24600
rect -386 -25052 302 -24628
rect 366 -25052 386 -24628
rect -386 -25080 386 -25052
rect -386 -25348 386 -25320
rect -386 -25772 302 -25348
rect 366 -25772 386 -25348
rect -386 -25800 386 -25772
rect -386 -26068 386 -26040
rect -386 -26492 302 -26068
rect 366 -26492 386 -26068
rect -386 -26520 386 -26492
rect -386 -26788 386 -26760
rect -386 -27212 302 -26788
rect 366 -27212 386 -26788
rect -386 -27240 386 -27212
rect -386 -27508 386 -27480
rect -386 -27932 302 -27508
rect 366 -27932 386 -27508
rect -386 -27960 386 -27932
rect -386 -28228 386 -28200
rect -386 -28652 302 -28228
rect 366 -28652 386 -28228
rect -386 -28680 386 -28652
rect -386 -28948 386 -28920
rect -386 -29372 302 -28948
rect 366 -29372 386 -28948
rect -386 -29400 386 -29372
rect -386 -29668 386 -29640
rect -386 -30092 302 -29668
rect 366 -30092 386 -29668
rect -386 -30120 386 -30092
rect -386 -30388 386 -30360
rect -386 -30812 302 -30388
rect 366 -30812 386 -30388
rect -386 -30840 386 -30812
rect -386 -31108 386 -31080
rect -386 -31532 302 -31108
rect 366 -31532 386 -31108
rect -386 -31560 386 -31532
rect -386 -31828 386 -31800
rect -386 -32252 302 -31828
rect 366 -32252 386 -31828
rect -386 -32280 386 -32252
rect -386 -32548 386 -32520
rect -386 -32972 302 -32548
rect 366 -32972 386 -32548
rect -386 -33000 386 -32972
rect -386 -33268 386 -33240
rect -386 -33692 302 -33268
rect 366 -33692 386 -33268
rect -386 -33720 386 -33692
rect -386 -33988 386 -33960
rect -386 -34412 302 -33988
rect 366 -34412 386 -33988
rect -386 -34440 386 -34412
rect -386 -34708 386 -34680
rect -386 -35132 302 -34708
rect 366 -35132 386 -34708
rect -386 -35160 386 -35132
rect -386 -35428 386 -35400
rect -386 -35852 302 -35428
rect 366 -35852 386 -35428
rect -386 -35880 386 -35852
rect -386 -36148 386 -36120
rect -386 -36572 302 -36148
rect 366 -36572 386 -36148
rect -386 -36600 386 -36572
rect -386 -36868 386 -36840
rect -386 -37292 302 -36868
rect 366 -37292 386 -36868
rect -386 -37320 386 -37292
rect -386 -37588 386 -37560
rect -386 -38012 302 -37588
rect 366 -38012 386 -37588
rect -386 -38040 386 -38012
rect -386 -38308 386 -38280
rect -386 -38732 302 -38308
rect 366 -38732 386 -38308
rect -386 -38760 386 -38732
rect -386 -39028 386 -39000
rect -386 -39452 302 -39028
rect 366 -39452 386 -39028
rect -386 -39480 386 -39452
rect -386 -39748 386 -39720
rect -386 -40172 302 -39748
rect 366 -40172 386 -39748
rect -386 -40200 386 -40172
rect -386 -40468 386 -40440
rect -386 -40892 302 -40468
rect 366 -40892 386 -40468
rect -386 -40920 386 -40892
rect -386 -41188 386 -41160
rect -386 -41612 302 -41188
rect 366 -41612 386 -41188
rect -386 -41640 386 -41612
rect -386 -41908 386 -41880
rect -386 -42332 302 -41908
rect 366 -42332 386 -41908
rect -386 -42360 386 -42332
rect -386 -42628 386 -42600
rect -386 -43052 302 -42628
rect 366 -43052 386 -42628
rect -386 -43080 386 -43052
rect -386 -43348 386 -43320
rect -386 -43772 302 -43348
rect 366 -43772 386 -43348
rect -386 -43800 386 -43772
rect -386 -44068 386 -44040
rect -386 -44492 302 -44068
rect 366 -44492 386 -44068
rect -386 -44520 386 -44492
rect -386 -44788 386 -44760
rect -386 -45212 302 -44788
rect 366 -45212 386 -44788
rect -386 -45240 386 -45212
rect -386 -45508 386 -45480
rect -386 -45932 302 -45508
rect 366 -45932 386 -45508
rect -386 -45960 386 -45932
<< via3 >>
rect 302 45508 366 45932
rect 302 44788 366 45212
rect 302 44068 366 44492
rect 302 43348 366 43772
rect 302 42628 366 43052
rect 302 41908 366 42332
rect 302 41188 366 41612
rect 302 40468 366 40892
rect 302 39748 366 40172
rect 302 39028 366 39452
rect 302 38308 366 38732
rect 302 37588 366 38012
rect 302 36868 366 37292
rect 302 36148 366 36572
rect 302 35428 366 35852
rect 302 34708 366 35132
rect 302 33988 366 34412
rect 302 33268 366 33692
rect 302 32548 366 32972
rect 302 31828 366 32252
rect 302 31108 366 31532
rect 302 30388 366 30812
rect 302 29668 366 30092
rect 302 28948 366 29372
rect 302 28228 366 28652
rect 302 27508 366 27932
rect 302 26788 366 27212
rect 302 26068 366 26492
rect 302 25348 366 25772
rect 302 24628 366 25052
rect 302 23908 366 24332
rect 302 23188 366 23612
rect 302 22468 366 22892
rect 302 21748 366 22172
rect 302 21028 366 21452
rect 302 20308 366 20732
rect 302 19588 366 20012
rect 302 18868 366 19292
rect 302 18148 366 18572
rect 302 17428 366 17852
rect 302 16708 366 17132
rect 302 15988 366 16412
rect 302 15268 366 15692
rect 302 14548 366 14972
rect 302 13828 366 14252
rect 302 13108 366 13532
rect 302 12388 366 12812
rect 302 11668 366 12092
rect 302 10948 366 11372
rect 302 10228 366 10652
rect 302 9508 366 9932
rect 302 8788 366 9212
rect 302 8068 366 8492
rect 302 7348 366 7772
rect 302 6628 366 7052
rect 302 5908 366 6332
rect 302 5188 366 5612
rect 302 4468 366 4892
rect 302 3748 366 4172
rect 302 3028 366 3452
rect 302 2308 366 2732
rect 302 1588 366 2012
rect 302 868 366 1292
rect 302 148 366 572
rect 302 -572 366 -148
rect 302 -1292 366 -868
rect 302 -2012 366 -1588
rect 302 -2732 366 -2308
rect 302 -3452 366 -3028
rect 302 -4172 366 -3748
rect 302 -4892 366 -4468
rect 302 -5612 366 -5188
rect 302 -6332 366 -5908
rect 302 -7052 366 -6628
rect 302 -7772 366 -7348
rect 302 -8492 366 -8068
rect 302 -9212 366 -8788
rect 302 -9932 366 -9508
rect 302 -10652 366 -10228
rect 302 -11372 366 -10948
rect 302 -12092 366 -11668
rect 302 -12812 366 -12388
rect 302 -13532 366 -13108
rect 302 -14252 366 -13828
rect 302 -14972 366 -14548
rect 302 -15692 366 -15268
rect 302 -16412 366 -15988
rect 302 -17132 366 -16708
rect 302 -17852 366 -17428
rect 302 -18572 366 -18148
rect 302 -19292 366 -18868
rect 302 -20012 366 -19588
rect 302 -20732 366 -20308
rect 302 -21452 366 -21028
rect 302 -22172 366 -21748
rect 302 -22892 366 -22468
rect 302 -23612 366 -23188
rect 302 -24332 366 -23908
rect 302 -25052 366 -24628
rect 302 -25772 366 -25348
rect 302 -26492 366 -26068
rect 302 -27212 366 -26788
rect 302 -27932 366 -27508
rect 302 -28652 366 -28228
rect 302 -29372 366 -28948
rect 302 -30092 366 -29668
rect 302 -30812 366 -30388
rect 302 -31532 366 -31108
rect 302 -32252 366 -31828
rect 302 -32972 366 -32548
rect 302 -33692 366 -33268
rect 302 -34412 366 -33988
rect 302 -35132 366 -34708
rect 302 -35852 366 -35428
rect 302 -36572 366 -36148
rect 302 -37292 366 -36868
rect 302 -38012 366 -37588
rect 302 -38732 366 -38308
rect 302 -39452 366 -39028
rect 302 -40172 366 -39748
rect 302 -40892 366 -40468
rect 302 -41612 366 -41188
rect 302 -42332 366 -41908
rect 302 -43052 366 -42628
rect 302 -43772 366 -43348
rect 302 -44492 366 -44068
rect 302 -45212 366 -44788
rect 302 -45932 366 -45508
<< mimcap >>
rect -346 45880 54 45920
rect -346 45560 -306 45880
rect 14 45560 54 45880
rect -346 45520 54 45560
rect -346 45160 54 45200
rect -346 44840 -306 45160
rect 14 44840 54 45160
rect -346 44800 54 44840
rect -346 44440 54 44480
rect -346 44120 -306 44440
rect 14 44120 54 44440
rect -346 44080 54 44120
rect -346 43720 54 43760
rect -346 43400 -306 43720
rect 14 43400 54 43720
rect -346 43360 54 43400
rect -346 43000 54 43040
rect -346 42680 -306 43000
rect 14 42680 54 43000
rect -346 42640 54 42680
rect -346 42280 54 42320
rect -346 41960 -306 42280
rect 14 41960 54 42280
rect -346 41920 54 41960
rect -346 41560 54 41600
rect -346 41240 -306 41560
rect 14 41240 54 41560
rect -346 41200 54 41240
rect -346 40840 54 40880
rect -346 40520 -306 40840
rect 14 40520 54 40840
rect -346 40480 54 40520
rect -346 40120 54 40160
rect -346 39800 -306 40120
rect 14 39800 54 40120
rect -346 39760 54 39800
rect -346 39400 54 39440
rect -346 39080 -306 39400
rect 14 39080 54 39400
rect -346 39040 54 39080
rect -346 38680 54 38720
rect -346 38360 -306 38680
rect 14 38360 54 38680
rect -346 38320 54 38360
rect -346 37960 54 38000
rect -346 37640 -306 37960
rect 14 37640 54 37960
rect -346 37600 54 37640
rect -346 37240 54 37280
rect -346 36920 -306 37240
rect 14 36920 54 37240
rect -346 36880 54 36920
rect -346 36520 54 36560
rect -346 36200 -306 36520
rect 14 36200 54 36520
rect -346 36160 54 36200
rect -346 35800 54 35840
rect -346 35480 -306 35800
rect 14 35480 54 35800
rect -346 35440 54 35480
rect -346 35080 54 35120
rect -346 34760 -306 35080
rect 14 34760 54 35080
rect -346 34720 54 34760
rect -346 34360 54 34400
rect -346 34040 -306 34360
rect 14 34040 54 34360
rect -346 34000 54 34040
rect -346 33640 54 33680
rect -346 33320 -306 33640
rect 14 33320 54 33640
rect -346 33280 54 33320
rect -346 32920 54 32960
rect -346 32600 -306 32920
rect 14 32600 54 32920
rect -346 32560 54 32600
rect -346 32200 54 32240
rect -346 31880 -306 32200
rect 14 31880 54 32200
rect -346 31840 54 31880
rect -346 31480 54 31520
rect -346 31160 -306 31480
rect 14 31160 54 31480
rect -346 31120 54 31160
rect -346 30760 54 30800
rect -346 30440 -306 30760
rect 14 30440 54 30760
rect -346 30400 54 30440
rect -346 30040 54 30080
rect -346 29720 -306 30040
rect 14 29720 54 30040
rect -346 29680 54 29720
rect -346 29320 54 29360
rect -346 29000 -306 29320
rect 14 29000 54 29320
rect -346 28960 54 29000
rect -346 28600 54 28640
rect -346 28280 -306 28600
rect 14 28280 54 28600
rect -346 28240 54 28280
rect -346 27880 54 27920
rect -346 27560 -306 27880
rect 14 27560 54 27880
rect -346 27520 54 27560
rect -346 27160 54 27200
rect -346 26840 -306 27160
rect 14 26840 54 27160
rect -346 26800 54 26840
rect -346 26440 54 26480
rect -346 26120 -306 26440
rect 14 26120 54 26440
rect -346 26080 54 26120
rect -346 25720 54 25760
rect -346 25400 -306 25720
rect 14 25400 54 25720
rect -346 25360 54 25400
rect -346 25000 54 25040
rect -346 24680 -306 25000
rect 14 24680 54 25000
rect -346 24640 54 24680
rect -346 24280 54 24320
rect -346 23960 -306 24280
rect 14 23960 54 24280
rect -346 23920 54 23960
rect -346 23560 54 23600
rect -346 23240 -306 23560
rect 14 23240 54 23560
rect -346 23200 54 23240
rect -346 22840 54 22880
rect -346 22520 -306 22840
rect 14 22520 54 22840
rect -346 22480 54 22520
rect -346 22120 54 22160
rect -346 21800 -306 22120
rect 14 21800 54 22120
rect -346 21760 54 21800
rect -346 21400 54 21440
rect -346 21080 -306 21400
rect 14 21080 54 21400
rect -346 21040 54 21080
rect -346 20680 54 20720
rect -346 20360 -306 20680
rect 14 20360 54 20680
rect -346 20320 54 20360
rect -346 19960 54 20000
rect -346 19640 -306 19960
rect 14 19640 54 19960
rect -346 19600 54 19640
rect -346 19240 54 19280
rect -346 18920 -306 19240
rect 14 18920 54 19240
rect -346 18880 54 18920
rect -346 18520 54 18560
rect -346 18200 -306 18520
rect 14 18200 54 18520
rect -346 18160 54 18200
rect -346 17800 54 17840
rect -346 17480 -306 17800
rect 14 17480 54 17800
rect -346 17440 54 17480
rect -346 17080 54 17120
rect -346 16760 -306 17080
rect 14 16760 54 17080
rect -346 16720 54 16760
rect -346 16360 54 16400
rect -346 16040 -306 16360
rect 14 16040 54 16360
rect -346 16000 54 16040
rect -346 15640 54 15680
rect -346 15320 -306 15640
rect 14 15320 54 15640
rect -346 15280 54 15320
rect -346 14920 54 14960
rect -346 14600 -306 14920
rect 14 14600 54 14920
rect -346 14560 54 14600
rect -346 14200 54 14240
rect -346 13880 -306 14200
rect 14 13880 54 14200
rect -346 13840 54 13880
rect -346 13480 54 13520
rect -346 13160 -306 13480
rect 14 13160 54 13480
rect -346 13120 54 13160
rect -346 12760 54 12800
rect -346 12440 -306 12760
rect 14 12440 54 12760
rect -346 12400 54 12440
rect -346 12040 54 12080
rect -346 11720 -306 12040
rect 14 11720 54 12040
rect -346 11680 54 11720
rect -346 11320 54 11360
rect -346 11000 -306 11320
rect 14 11000 54 11320
rect -346 10960 54 11000
rect -346 10600 54 10640
rect -346 10280 -306 10600
rect 14 10280 54 10600
rect -346 10240 54 10280
rect -346 9880 54 9920
rect -346 9560 -306 9880
rect 14 9560 54 9880
rect -346 9520 54 9560
rect -346 9160 54 9200
rect -346 8840 -306 9160
rect 14 8840 54 9160
rect -346 8800 54 8840
rect -346 8440 54 8480
rect -346 8120 -306 8440
rect 14 8120 54 8440
rect -346 8080 54 8120
rect -346 7720 54 7760
rect -346 7400 -306 7720
rect 14 7400 54 7720
rect -346 7360 54 7400
rect -346 7000 54 7040
rect -346 6680 -306 7000
rect 14 6680 54 7000
rect -346 6640 54 6680
rect -346 6280 54 6320
rect -346 5960 -306 6280
rect 14 5960 54 6280
rect -346 5920 54 5960
rect -346 5560 54 5600
rect -346 5240 -306 5560
rect 14 5240 54 5560
rect -346 5200 54 5240
rect -346 4840 54 4880
rect -346 4520 -306 4840
rect 14 4520 54 4840
rect -346 4480 54 4520
rect -346 4120 54 4160
rect -346 3800 -306 4120
rect 14 3800 54 4120
rect -346 3760 54 3800
rect -346 3400 54 3440
rect -346 3080 -306 3400
rect 14 3080 54 3400
rect -346 3040 54 3080
rect -346 2680 54 2720
rect -346 2360 -306 2680
rect 14 2360 54 2680
rect -346 2320 54 2360
rect -346 1960 54 2000
rect -346 1640 -306 1960
rect 14 1640 54 1960
rect -346 1600 54 1640
rect -346 1240 54 1280
rect -346 920 -306 1240
rect 14 920 54 1240
rect -346 880 54 920
rect -346 520 54 560
rect -346 200 -306 520
rect 14 200 54 520
rect -346 160 54 200
rect -346 -200 54 -160
rect -346 -520 -306 -200
rect 14 -520 54 -200
rect -346 -560 54 -520
rect -346 -920 54 -880
rect -346 -1240 -306 -920
rect 14 -1240 54 -920
rect -346 -1280 54 -1240
rect -346 -1640 54 -1600
rect -346 -1960 -306 -1640
rect 14 -1960 54 -1640
rect -346 -2000 54 -1960
rect -346 -2360 54 -2320
rect -346 -2680 -306 -2360
rect 14 -2680 54 -2360
rect -346 -2720 54 -2680
rect -346 -3080 54 -3040
rect -346 -3400 -306 -3080
rect 14 -3400 54 -3080
rect -346 -3440 54 -3400
rect -346 -3800 54 -3760
rect -346 -4120 -306 -3800
rect 14 -4120 54 -3800
rect -346 -4160 54 -4120
rect -346 -4520 54 -4480
rect -346 -4840 -306 -4520
rect 14 -4840 54 -4520
rect -346 -4880 54 -4840
rect -346 -5240 54 -5200
rect -346 -5560 -306 -5240
rect 14 -5560 54 -5240
rect -346 -5600 54 -5560
rect -346 -5960 54 -5920
rect -346 -6280 -306 -5960
rect 14 -6280 54 -5960
rect -346 -6320 54 -6280
rect -346 -6680 54 -6640
rect -346 -7000 -306 -6680
rect 14 -7000 54 -6680
rect -346 -7040 54 -7000
rect -346 -7400 54 -7360
rect -346 -7720 -306 -7400
rect 14 -7720 54 -7400
rect -346 -7760 54 -7720
rect -346 -8120 54 -8080
rect -346 -8440 -306 -8120
rect 14 -8440 54 -8120
rect -346 -8480 54 -8440
rect -346 -8840 54 -8800
rect -346 -9160 -306 -8840
rect 14 -9160 54 -8840
rect -346 -9200 54 -9160
rect -346 -9560 54 -9520
rect -346 -9880 -306 -9560
rect 14 -9880 54 -9560
rect -346 -9920 54 -9880
rect -346 -10280 54 -10240
rect -346 -10600 -306 -10280
rect 14 -10600 54 -10280
rect -346 -10640 54 -10600
rect -346 -11000 54 -10960
rect -346 -11320 -306 -11000
rect 14 -11320 54 -11000
rect -346 -11360 54 -11320
rect -346 -11720 54 -11680
rect -346 -12040 -306 -11720
rect 14 -12040 54 -11720
rect -346 -12080 54 -12040
rect -346 -12440 54 -12400
rect -346 -12760 -306 -12440
rect 14 -12760 54 -12440
rect -346 -12800 54 -12760
rect -346 -13160 54 -13120
rect -346 -13480 -306 -13160
rect 14 -13480 54 -13160
rect -346 -13520 54 -13480
rect -346 -13880 54 -13840
rect -346 -14200 -306 -13880
rect 14 -14200 54 -13880
rect -346 -14240 54 -14200
rect -346 -14600 54 -14560
rect -346 -14920 -306 -14600
rect 14 -14920 54 -14600
rect -346 -14960 54 -14920
rect -346 -15320 54 -15280
rect -346 -15640 -306 -15320
rect 14 -15640 54 -15320
rect -346 -15680 54 -15640
rect -346 -16040 54 -16000
rect -346 -16360 -306 -16040
rect 14 -16360 54 -16040
rect -346 -16400 54 -16360
rect -346 -16760 54 -16720
rect -346 -17080 -306 -16760
rect 14 -17080 54 -16760
rect -346 -17120 54 -17080
rect -346 -17480 54 -17440
rect -346 -17800 -306 -17480
rect 14 -17800 54 -17480
rect -346 -17840 54 -17800
rect -346 -18200 54 -18160
rect -346 -18520 -306 -18200
rect 14 -18520 54 -18200
rect -346 -18560 54 -18520
rect -346 -18920 54 -18880
rect -346 -19240 -306 -18920
rect 14 -19240 54 -18920
rect -346 -19280 54 -19240
rect -346 -19640 54 -19600
rect -346 -19960 -306 -19640
rect 14 -19960 54 -19640
rect -346 -20000 54 -19960
rect -346 -20360 54 -20320
rect -346 -20680 -306 -20360
rect 14 -20680 54 -20360
rect -346 -20720 54 -20680
rect -346 -21080 54 -21040
rect -346 -21400 -306 -21080
rect 14 -21400 54 -21080
rect -346 -21440 54 -21400
rect -346 -21800 54 -21760
rect -346 -22120 -306 -21800
rect 14 -22120 54 -21800
rect -346 -22160 54 -22120
rect -346 -22520 54 -22480
rect -346 -22840 -306 -22520
rect 14 -22840 54 -22520
rect -346 -22880 54 -22840
rect -346 -23240 54 -23200
rect -346 -23560 -306 -23240
rect 14 -23560 54 -23240
rect -346 -23600 54 -23560
rect -346 -23960 54 -23920
rect -346 -24280 -306 -23960
rect 14 -24280 54 -23960
rect -346 -24320 54 -24280
rect -346 -24680 54 -24640
rect -346 -25000 -306 -24680
rect 14 -25000 54 -24680
rect -346 -25040 54 -25000
rect -346 -25400 54 -25360
rect -346 -25720 -306 -25400
rect 14 -25720 54 -25400
rect -346 -25760 54 -25720
rect -346 -26120 54 -26080
rect -346 -26440 -306 -26120
rect 14 -26440 54 -26120
rect -346 -26480 54 -26440
rect -346 -26840 54 -26800
rect -346 -27160 -306 -26840
rect 14 -27160 54 -26840
rect -346 -27200 54 -27160
rect -346 -27560 54 -27520
rect -346 -27880 -306 -27560
rect 14 -27880 54 -27560
rect -346 -27920 54 -27880
rect -346 -28280 54 -28240
rect -346 -28600 -306 -28280
rect 14 -28600 54 -28280
rect -346 -28640 54 -28600
rect -346 -29000 54 -28960
rect -346 -29320 -306 -29000
rect 14 -29320 54 -29000
rect -346 -29360 54 -29320
rect -346 -29720 54 -29680
rect -346 -30040 -306 -29720
rect 14 -30040 54 -29720
rect -346 -30080 54 -30040
rect -346 -30440 54 -30400
rect -346 -30760 -306 -30440
rect 14 -30760 54 -30440
rect -346 -30800 54 -30760
rect -346 -31160 54 -31120
rect -346 -31480 -306 -31160
rect 14 -31480 54 -31160
rect -346 -31520 54 -31480
rect -346 -31880 54 -31840
rect -346 -32200 -306 -31880
rect 14 -32200 54 -31880
rect -346 -32240 54 -32200
rect -346 -32600 54 -32560
rect -346 -32920 -306 -32600
rect 14 -32920 54 -32600
rect -346 -32960 54 -32920
rect -346 -33320 54 -33280
rect -346 -33640 -306 -33320
rect 14 -33640 54 -33320
rect -346 -33680 54 -33640
rect -346 -34040 54 -34000
rect -346 -34360 -306 -34040
rect 14 -34360 54 -34040
rect -346 -34400 54 -34360
rect -346 -34760 54 -34720
rect -346 -35080 -306 -34760
rect 14 -35080 54 -34760
rect -346 -35120 54 -35080
rect -346 -35480 54 -35440
rect -346 -35800 -306 -35480
rect 14 -35800 54 -35480
rect -346 -35840 54 -35800
rect -346 -36200 54 -36160
rect -346 -36520 -306 -36200
rect 14 -36520 54 -36200
rect -346 -36560 54 -36520
rect -346 -36920 54 -36880
rect -346 -37240 -306 -36920
rect 14 -37240 54 -36920
rect -346 -37280 54 -37240
rect -346 -37640 54 -37600
rect -346 -37960 -306 -37640
rect 14 -37960 54 -37640
rect -346 -38000 54 -37960
rect -346 -38360 54 -38320
rect -346 -38680 -306 -38360
rect 14 -38680 54 -38360
rect -346 -38720 54 -38680
rect -346 -39080 54 -39040
rect -346 -39400 -306 -39080
rect 14 -39400 54 -39080
rect -346 -39440 54 -39400
rect -346 -39800 54 -39760
rect -346 -40120 -306 -39800
rect 14 -40120 54 -39800
rect -346 -40160 54 -40120
rect -346 -40520 54 -40480
rect -346 -40840 -306 -40520
rect 14 -40840 54 -40520
rect -346 -40880 54 -40840
rect -346 -41240 54 -41200
rect -346 -41560 -306 -41240
rect 14 -41560 54 -41240
rect -346 -41600 54 -41560
rect -346 -41960 54 -41920
rect -346 -42280 -306 -41960
rect 14 -42280 54 -41960
rect -346 -42320 54 -42280
rect -346 -42680 54 -42640
rect -346 -43000 -306 -42680
rect 14 -43000 54 -42680
rect -346 -43040 54 -43000
rect -346 -43400 54 -43360
rect -346 -43720 -306 -43400
rect 14 -43720 54 -43400
rect -346 -43760 54 -43720
rect -346 -44120 54 -44080
rect -346 -44440 -306 -44120
rect 14 -44440 54 -44120
rect -346 -44480 54 -44440
rect -346 -44840 54 -44800
rect -346 -45160 -306 -44840
rect 14 -45160 54 -44840
rect -346 -45200 54 -45160
rect -346 -45560 54 -45520
rect -346 -45880 -306 -45560
rect 14 -45880 54 -45560
rect -346 -45920 54 -45880
<< mimcapcontact >>
rect -306 45560 14 45880
rect -306 44840 14 45160
rect -306 44120 14 44440
rect -306 43400 14 43720
rect -306 42680 14 43000
rect -306 41960 14 42280
rect -306 41240 14 41560
rect -306 40520 14 40840
rect -306 39800 14 40120
rect -306 39080 14 39400
rect -306 38360 14 38680
rect -306 37640 14 37960
rect -306 36920 14 37240
rect -306 36200 14 36520
rect -306 35480 14 35800
rect -306 34760 14 35080
rect -306 34040 14 34360
rect -306 33320 14 33640
rect -306 32600 14 32920
rect -306 31880 14 32200
rect -306 31160 14 31480
rect -306 30440 14 30760
rect -306 29720 14 30040
rect -306 29000 14 29320
rect -306 28280 14 28600
rect -306 27560 14 27880
rect -306 26840 14 27160
rect -306 26120 14 26440
rect -306 25400 14 25720
rect -306 24680 14 25000
rect -306 23960 14 24280
rect -306 23240 14 23560
rect -306 22520 14 22840
rect -306 21800 14 22120
rect -306 21080 14 21400
rect -306 20360 14 20680
rect -306 19640 14 19960
rect -306 18920 14 19240
rect -306 18200 14 18520
rect -306 17480 14 17800
rect -306 16760 14 17080
rect -306 16040 14 16360
rect -306 15320 14 15640
rect -306 14600 14 14920
rect -306 13880 14 14200
rect -306 13160 14 13480
rect -306 12440 14 12760
rect -306 11720 14 12040
rect -306 11000 14 11320
rect -306 10280 14 10600
rect -306 9560 14 9880
rect -306 8840 14 9160
rect -306 8120 14 8440
rect -306 7400 14 7720
rect -306 6680 14 7000
rect -306 5960 14 6280
rect -306 5240 14 5560
rect -306 4520 14 4840
rect -306 3800 14 4120
rect -306 3080 14 3400
rect -306 2360 14 2680
rect -306 1640 14 1960
rect -306 920 14 1240
rect -306 200 14 520
rect -306 -520 14 -200
rect -306 -1240 14 -920
rect -306 -1960 14 -1640
rect -306 -2680 14 -2360
rect -306 -3400 14 -3080
rect -306 -4120 14 -3800
rect -306 -4840 14 -4520
rect -306 -5560 14 -5240
rect -306 -6280 14 -5960
rect -306 -7000 14 -6680
rect -306 -7720 14 -7400
rect -306 -8440 14 -8120
rect -306 -9160 14 -8840
rect -306 -9880 14 -9560
rect -306 -10600 14 -10280
rect -306 -11320 14 -11000
rect -306 -12040 14 -11720
rect -306 -12760 14 -12440
rect -306 -13480 14 -13160
rect -306 -14200 14 -13880
rect -306 -14920 14 -14600
rect -306 -15640 14 -15320
rect -306 -16360 14 -16040
rect -306 -17080 14 -16760
rect -306 -17800 14 -17480
rect -306 -18520 14 -18200
rect -306 -19240 14 -18920
rect -306 -19960 14 -19640
rect -306 -20680 14 -20360
rect -306 -21400 14 -21080
rect -306 -22120 14 -21800
rect -306 -22840 14 -22520
rect -306 -23560 14 -23240
rect -306 -24280 14 -23960
rect -306 -25000 14 -24680
rect -306 -25720 14 -25400
rect -306 -26440 14 -26120
rect -306 -27160 14 -26840
rect -306 -27880 14 -27560
rect -306 -28600 14 -28280
rect -306 -29320 14 -29000
rect -306 -30040 14 -29720
rect -306 -30760 14 -30440
rect -306 -31480 14 -31160
rect -306 -32200 14 -31880
rect -306 -32920 14 -32600
rect -306 -33640 14 -33320
rect -306 -34360 14 -34040
rect -306 -35080 14 -34760
rect -306 -35800 14 -35480
rect -306 -36520 14 -36200
rect -306 -37240 14 -36920
rect -306 -37960 14 -37640
rect -306 -38680 14 -38360
rect -306 -39400 14 -39080
rect -306 -40120 14 -39800
rect -306 -40840 14 -40520
rect -306 -41560 14 -41240
rect -306 -42280 14 -41960
rect -306 -43000 14 -42680
rect -306 -43720 14 -43400
rect -306 -44440 14 -44120
rect -306 -45160 14 -44840
rect -306 -45880 14 -45560
<< metal4 >>
rect -198 45881 -94 46080
rect 282 45932 386 46080
rect -307 45880 15 45881
rect -307 45560 -306 45880
rect 14 45560 15 45880
rect -307 45559 15 45560
rect -198 45161 -94 45559
rect 282 45508 302 45932
rect 366 45508 386 45932
rect 282 45212 386 45508
rect -307 45160 15 45161
rect -307 44840 -306 45160
rect 14 44840 15 45160
rect -307 44839 15 44840
rect -198 44441 -94 44839
rect 282 44788 302 45212
rect 366 44788 386 45212
rect 282 44492 386 44788
rect -307 44440 15 44441
rect -307 44120 -306 44440
rect 14 44120 15 44440
rect -307 44119 15 44120
rect -198 43721 -94 44119
rect 282 44068 302 44492
rect 366 44068 386 44492
rect 282 43772 386 44068
rect -307 43720 15 43721
rect -307 43400 -306 43720
rect 14 43400 15 43720
rect -307 43399 15 43400
rect -198 43001 -94 43399
rect 282 43348 302 43772
rect 366 43348 386 43772
rect 282 43052 386 43348
rect -307 43000 15 43001
rect -307 42680 -306 43000
rect 14 42680 15 43000
rect -307 42679 15 42680
rect -198 42281 -94 42679
rect 282 42628 302 43052
rect 366 42628 386 43052
rect 282 42332 386 42628
rect -307 42280 15 42281
rect -307 41960 -306 42280
rect 14 41960 15 42280
rect -307 41959 15 41960
rect -198 41561 -94 41959
rect 282 41908 302 42332
rect 366 41908 386 42332
rect 282 41612 386 41908
rect -307 41560 15 41561
rect -307 41240 -306 41560
rect 14 41240 15 41560
rect -307 41239 15 41240
rect -198 40841 -94 41239
rect 282 41188 302 41612
rect 366 41188 386 41612
rect 282 40892 386 41188
rect -307 40840 15 40841
rect -307 40520 -306 40840
rect 14 40520 15 40840
rect -307 40519 15 40520
rect -198 40121 -94 40519
rect 282 40468 302 40892
rect 366 40468 386 40892
rect 282 40172 386 40468
rect -307 40120 15 40121
rect -307 39800 -306 40120
rect 14 39800 15 40120
rect -307 39799 15 39800
rect -198 39401 -94 39799
rect 282 39748 302 40172
rect 366 39748 386 40172
rect 282 39452 386 39748
rect -307 39400 15 39401
rect -307 39080 -306 39400
rect 14 39080 15 39400
rect -307 39079 15 39080
rect -198 38681 -94 39079
rect 282 39028 302 39452
rect 366 39028 386 39452
rect 282 38732 386 39028
rect -307 38680 15 38681
rect -307 38360 -306 38680
rect 14 38360 15 38680
rect -307 38359 15 38360
rect -198 37961 -94 38359
rect 282 38308 302 38732
rect 366 38308 386 38732
rect 282 38012 386 38308
rect -307 37960 15 37961
rect -307 37640 -306 37960
rect 14 37640 15 37960
rect -307 37639 15 37640
rect -198 37241 -94 37639
rect 282 37588 302 38012
rect 366 37588 386 38012
rect 282 37292 386 37588
rect -307 37240 15 37241
rect -307 36920 -306 37240
rect 14 36920 15 37240
rect -307 36919 15 36920
rect -198 36521 -94 36919
rect 282 36868 302 37292
rect 366 36868 386 37292
rect 282 36572 386 36868
rect -307 36520 15 36521
rect -307 36200 -306 36520
rect 14 36200 15 36520
rect -307 36199 15 36200
rect -198 35801 -94 36199
rect 282 36148 302 36572
rect 366 36148 386 36572
rect 282 35852 386 36148
rect -307 35800 15 35801
rect -307 35480 -306 35800
rect 14 35480 15 35800
rect -307 35479 15 35480
rect -198 35081 -94 35479
rect 282 35428 302 35852
rect 366 35428 386 35852
rect 282 35132 386 35428
rect -307 35080 15 35081
rect -307 34760 -306 35080
rect 14 34760 15 35080
rect -307 34759 15 34760
rect -198 34361 -94 34759
rect 282 34708 302 35132
rect 366 34708 386 35132
rect 282 34412 386 34708
rect -307 34360 15 34361
rect -307 34040 -306 34360
rect 14 34040 15 34360
rect -307 34039 15 34040
rect -198 33641 -94 34039
rect 282 33988 302 34412
rect 366 33988 386 34412
rect 282 33692 386 33988
rect -307 33640 15 33641
rect -307 33320 -306 33640
rect 14 33320 15 33640
rect -307 33319 15 33320
rect -198 32921 -94 33319
rect 282 33268 302 33692
rect 366 33268 386 33692
rect 282 32972 386 33268
rect -307 32920 15 32921
rect -307 32600 -306 32920
rect 14 32600 15 32920
rect -307 32599 15 32600
rect -198 32201 -94 32599
rect 282 32548 302 32972
rect 366 32548 386 32972
rect 282 32252 386 32548
rect -307 32200 15 32201
rect -307 31880 -306 32200
rect 14 31880 15 32200
rect -307 31879 15 31880
rect -198 31481 -94 31879
rect 282 31828 302 32252
rect 366 31828 386 32252
rect 282 31532 386 31828
rect -307 31480 15 31481
rect -307 31160 -306 31480
rect 14 31160 15 31480
rect -307 31159 15 31160
rect -198 30761 -94 31159
rect 282 31108 302 31532
rect 366 31108 386 31532
rect 282 30812 386 31108
rect -307 30760 15 30761
rect -307 30440 -306 30760
rect 14 30440 15 30760
rect -307 30439 15 30440
rect -198 30041 -94 30439
rect 282 30388 302 30812
rect 366 30388 386 30812
rect 282 30092 386 30388
rect -307 30040 15 30041
rect -307 29720 -306 30040
rect 14 29720 15 30040
rect -307 29719 15 29720
rect -198 29321 -94 29719
rect 282 29668 302 30092
rect 366 29668 386 30092
rect 282 29372 386 29668
rect -307 29320 15 29321
rect -307 29000 -306 29320
rect 14 29000 15 29320
rect -307 28999 15 29000
rect -198 28601 -94 28999
rect 282 28948 302 29372
rect 366 28948 386 29372
rect 282 28652 386 28948
rect -307 28600 15 28601
rect -307 28280 -306 28600
rect 14 28280 15 28600
rect -307 28279 15 28280
rect -198 27881 -94 28279
rect 282 28228 302 28652
rect 366 28228 386 28652
rect 282 27932 386 28228
rect -307 27880 15 27881
rect -307 27560 -306 27880
rect 14 27560 15 27880
rect -307 27559 15 27560
rect -198 27161 -94 27559
rect 282 27508 302 27932
rect 366 27508 386 27932
rect 282 27212 386 27508
rect -307 27160 15 27161
rect -307 26840 -306 27160
rect 14 26840 15 27160
rect -307 26839 15 26840
rect -198 26441 -94 26839
rect 282 26788 302 27212
rect 366 26788 386 27212
rect 282 26492 386 26788
rect -307 26440 15 26441
rect -307 26120 -306 26440
rect 14 26120 15 26440
rect -307 26119 15 26120
rect -198 25721 -94 26119
rect 282 26068 302 26492
rect 366 26068 386 26492
rect 282 25772 386 26068
rect -307 25720 15 25721
rect -307 25400 -306 25720
rect 14 25400 15 25720
rect -307 25399 15 25400
rect -198 25001 -94 25399
rect 282 25348 302 25772
rect 366 25348 386 25772
rect 282 25052 386 25348
rect -307 25000 15 25001
rect -307 24680 -306 25000
rect 14 24680 15 25000
rect -307 24679 15 24680
rect -198 24281 -94 24679
rect 282 24628 302 25052
rect 366 24628 386 25052
rect 282 24332 386 24628
rect -307 24280 15 24281
rect -307 23960 -306 24280
rect 14 23960 15 24280
rect -307 23959 15 23960
rect -198 23561 -94 23959
rect 282 23908 302 24332
rect 366 23908 386 24332
rect 282 23612 386 23908
rect -307 23560 15 23561
rect -307 23240 -306 23560
rect 14 23240 15 23560
rect -307 23239 15 23240
rect -198 22841 -94 23239
rect 282 23188 302 23612
rect 366 23188 386 23612
rect 282 22892 386 23188
rect -307 22840 15 22841
rect -307 22520 -306 22840
rect 14 22520 15 22840
rect -307 22519 15 22520
rect -198 22121 -94 22519
rect 282 22468 302 22892
rect 366 22468 386 22892
rect 282 22172 386 22468
rect -307 22120 15 22121
rect -307 21800 -306 22120
rect 14 21800 15 22120
rect -307 21799 15 21800
rect -198 21401 -94 21799
rect 282 21748 302 22172
rect 366 21748 386 22172
rect 282 21452 386 21748
rect -307 21400 15 21401
rect -307 21080 -306 21400
rect 14 21080 15 21400
rect -307 21079 15 21080
rect -198 20681 -94 21079
rect 282 21028 302 21452
rect 366 21028 386 21452
rect 282 20732 386 21028
rect -307 20680 15 20681
rect -307 20360 -306 20680
rect 14 20360 15 20680
rect -307 20359 15 20360
rect -198 19961 -94 20359
rect 282 20308 302 20732
rect 366 20308 386 20732
rect 282 20012 386 20308
rect -307 19960 15 19961
rect -307 19640 -306 19960
rect 14 19640 15 19960
rect -307 19639 15 19640
rect -198 19241 -94 19639
rect 282 19588 302 20012
rect 366 19588 386 20012
rect 282 19292 386 19588
rect -307 19240 15 19241
rect -307 18920 -306 19240
rect 14 18920 15 19240
rect -307 18919 15 18920
rect -198 18521 -94 18919
rect 282 18868 302 19292
rect 366 18868 386 19292
rect 282 18572 386 18868
rect -307 18520 15 18521
rect -307 18200 -306 18520
rect 14 18200 15 18520
rect -307 18199 15 18200
rect -198 17801 -94 18199
rect 282 18148 302 18572
rect 366 18148 386 18572
rect 282 17852 386 18148
rect -307 17800 15 17801
rect -307 17480 -306 17800
rect 14 17480 15 17800
rect -307 17479 15 17480
rect -198 17081 -94 17479
rect 282 17428 302 17852
rect 366 17428 386 17852
rect 282 17132 386 17428
rect -307 17080 15 17081
rect -307 16760 -306 17080
rect 14 16760 15 17080
rect -307 16759 15 16760
rect -198 16361 -94 16759
rect 282 16708 302 17132
rect 366 16708 386 17132
rect 282 16412 386 16708
rect -307 16360 15 16361
rect -307 16040 -306 16360
rect 14 16040 15 16360
rect -307 16039 15 16040
rect -198 15641 -94 16039
rect 282 15988 302 16412
rect 366 15988 386 16412
rect 282 15692 386 15988
rect -307 15640 15 15641
rect -307 15320 -306 15640
rect 14 15320 15 15640
rect -307 15319 15 15320
rect -198 14921 -94 15319
rect 282 15268 302 15692
rect 366 15268 386 15692
rect 282 14972 386 15268
rect -307 14920 15 14921
rect -307 14600 -306 14920
rect 14 14600 15 14920
rect -307 14599 15 14600
rect -198 14201 -94 14599
rect 282 14548 302 14972
rect 366 14548 386 14972
rect 282 14252 386 14548
rect -307 14200 15 14201
rect -307 13880 -306 14200
rect 14 13880 15 14200
rect -307 13879 15 13880
rect -198 13481 -94 13879
rect 282 13828 302 14252
rect 366 13828 386 14252
rect 282 13532 386 13828
rect -307 13480 15 13481
rect -307 13160 -306 13480
rect 14 13160 15 13480
rect -307 13159 15 13160
rect -198 12761 -94 13159
rect 282 13108 302 13532
rect 366 13108 386 13532
rect 282 12812 386 13108
rect -307 12760 15 12761
rect -307 12440 -306 12760
rect 14 12440 15 12760
rect -307 12439 15 12440
rect -198 12041 -94 12439
rect 282 12388 302 12812
rect 366 12388 386 12812
rect 282 12092 386 12388
rect -307 12040 15 12041
rect -307 11720 -306 12040
rect 14 11720 15 12040
rect -307 11719 15 11720
rect -198 11321 -94 11719
rect 282 11668 302 12092
rect 366 11668 386 12092
rect 282 11372 386 11668
rect -307 11320 15 11321
rect -307 11000 -306 11320
rect 14 11000 15 11320
rect -307 10999 15 11000
rect -198 10601 -94 10999
rect 282 10948 302 11372
rect 366 10948 386 11372
rect 282 10652 386 10948
rect -307 10600 15 10601
rect -307 10280 -306 10600
rect 14 10280 15 10600
rect -307 10279 15 10280
rect -198 9881 -94 10279
rect 282 10228 302 10652
rect 366 10228 386 10652
rect 282 9932 386 10228
rect -307 9880 15 9881
rect -307 9560 -306 9880
rect 14 9560 15 9880
rect -307 9559 15 9560
rect -198 9161 -94 9559
rect 282 9508 302 9932
rect 366 9508 386 9932
rect 282 9212 386 9508
rect -307 9160 15 9161
rect -307 8840 -306 9160
rect 14 8840 15 9160
rect -307 8839 15 8840
rect -198 8441 -94 8839
rect 282 8788 302 9212
rect 366 8788 386 9212
rect 282 8492 386 8788
rect -307 8440 15 8441
rect -307 8120 -306 8440
rect 14 8120 15 8440
rect -307 8119 15 8120
rect -198 7721 -94 8119
rect 282 8068 302 8492
rect 366 8068 386 8492
rect 282 7772 386 8068
rect -307 7720 15 7721
rect -307 7400 -306 7720
rect 14 7400 15 7720
rect -307 7399 15 7400
rect -198 7001 -94 7399
rect 282 7348 302 7772
rect 366 7348 386 7772
rect 282 7052 386 7348
rect -307 7000 15 7001
rect -307 6680 -306 7000
rect 14 6680 15 7000
rect -307 6679 15 6680
rect -198 6281 -94 6679
rect 282 6628 302 7052
rect 366 6628 386 7052
rect 282 6332 386 6628
rect -307 6280 15 6281
rect -307 5960 -306 6280
rect 14 5960 15 6280
rect -307 5959 15 5960
rect -198 5561 -94 5959
rect 282 5908 302 6332
rect 366 5908 386 6332
rect 282 5612 386 5908
rect -307 5560 15 5561
rect -307 5240 -306 5560
rect 14 5240 15 5560
rect -307 5239 15 5240
rect -198 4841 -94 5239
rect 282 5188 302 5612
rect 366 5188 386 5612
rect 282 4892 386 5188
rect -307 4840 15 4841
rect -307 4520 -306 4840
rect 14 4520 15 4840
rect -307 4519 15 4520
rect -198 4121 -94 4519
rect 282 4468 302 4892
rect 366 4468 386 4892
rect 282 4172 386 4468
rect -307 4120 15 4121
rect -307 3800 -306 4120
rect 14 3800 15 4120
rect -307 3799 15 3800
rect -198 3401 -94 3799
rect 282 3748 302 4172
rect 366 3748 386 4172
rect 282 3452 386 3748
rect -307 3400 15 3401
rect -307 3080 -306 3400
rect 14 3080 15 3400
rect -307 3079 15 3080
rect -198 2681 -94 3079
rect 282 3028 302 3452
rect 366 3028 386 3452
rect 282 2732 386 3028
rect -307 2680 15 2681
rect -307 2360 -306 2680
rect 14 2360 15 2680
rect -307 2359 15 2360
rect -198 1961 -94 2359
rect 282 2308 302 2732
rect 366 2308 386 2732
rect 282 2012 386 2308
rect -307 1960 15 1961
rect -307 1640 -306 1960
rect 14 1640 15 1960
rect -307 1639 15 1640
rect -198 1241 -94 1639
rect 282 1588 302 2012
rect 366 1588 386 2012
rect 282 1292 386 1588
rect -307 1240 15 1241
rect -307 920 -306 1240
rect 14 920 15 1240
rect -307 919 15 920
rect -198 521 -94 919
rect 282 868 302 1292
rect 366 868 386 1292
rect 282 572 386 868
rect -307 520 15 521
rect -307 200 -306 520
rect 14 200 15 520
rect -307 199 15 200
rect -198 -199 -94 199
rect 282 148 302 572
rect 366 148 386 572
rect 282 -148 386 148
rect -307 -200 15 -199
rect -307 -520 -306 -200
rect 14 -520 15 -200
rect -307 -521 15 -520
rect -198 -919 -94 -521
rect 282 -572 302 -148
rect 366 -572 386 -148
rect 282 -868 386 -572
rect -307 -920 15 -919
rect -307 -1240 -306 -920
rect 14 -1240 15 -920
rect -307 -1241 15 -1240
rect -198 -1639 -94 -1241
rect 282 -1292 302 -868
rect 366 -1292 386 -868
rect 282 -1588 386 -1292
rect -307 -1640 15 -1639
rect -307 -1960 -306 -1640
rect 14 -1960 15 -1640
rect -307 -1961 15 -1960
rect -198 -2359 -94 -1961
rect 282 -2012 302 -1588
rect 366 -2012 386 -1588
rect 282 -2308 386 -2012
rect -307 -2360 15 -2359
rect -307 -2680 -306 -2360
rect 14 -2680 15 -2360
rect -307 -2681 15 -2680
rect -198 -3079 -94 -2681
rect 282 -2732 302 -2308
rect 366 -2732 386 -2308
rect 282 -3028 386 -2732
rect -307 -3080 15 -3079
rect -307 -3400 -306 -3080
rect 14 -3400 15 -3080
rect -307 -3401 15 -3400
rect -198 -3799 -94 -3401
rect 282 -3452 302 -3028
rect 366 -3452 386 -3028
rect 282 -3748 386 -3452
rect -307 -3800 15 -3799
rect -307 -4120 -306 -3800
rect 14 -4120 15 -3800
rect -307 -4121 15 -4120
rect -198 -4519 -94 -4121
rect 282 -4172 302 -3748
rect 366 -4172 386 -3748
rect 282 -4468 386 -4172
rect -307 -4520 15 -4519
rect -307 -4840 -306 -4520
rect 14 -4840 15 -4520
rect -307 -4841 15 -4840
rect -198 -5239 -94 -4841
rect 282 -4892 302 -4468
rect 366 -4892 386 -4468
rect 282 -5188 386 -4892
rect -307 -5240 15 -5239
rect -307 -5560 -306 -5240
rect 14 -5560 15 -5240
rect -307 -5561 15 -5560
rect -198 -5959 -94 -5561
rect 282 -5612 302 -5188
rect 366 -5612 386 -5188
rect 282 -5908 386 -5612
rect -307 -5960 15 -5959
rect -307 -6280 -306 -5960
rect 14 -6280 15 -5960
rect -307 -6281 15 -6280
rect -198 -6679 -94 -6281
rect 282 -6332 302 -5908
rect 366 -6332 386 -5908
rect 282 -6628 386 -6332
rect -307 -6680 15 -6679
rect -307 -7000 -306 -6680
rect 14 -7000 15 -6680
rect -307 -7001 15 -7000
rect -198 -7399 -94 -7001
rect 282 -7052 302 -6628
rect 366 -7052 386 -6628
rect 282 -7348 386 -7052
rect -307 -7400 15 -7399
rect -307 -7720 -306 -7400
rect 14 -7720 15 -7400
rect -307 -7721 15 -7720
rect -198 -8119 -94 -7721
rect 282 -7772 302 -7348
rect 366 -7772 386 -7348
rect 282 -8068 386 -7772
rect -307 -8120 15 -8119
rect -307 -8440 -306 -8120
rect 14 -8440 15 -8120
rect -307 -8441 15 -8440
rect -198 -8839 -94 -8441
rect 282 -8492 302 -8068
rect 366 -8492 386 -8068
rect 282 -8788 386 -8492
rect -307 -8840 15 -8839
rect -307 -9160 -306 -8840
rect 14 -9160 15 -8840
rect -307 -9161 15 -9160
rect -198 -9559 -94 -9161
rect 282 -9212 302 -8788
rect 366 -9212 386 -8788
rect 282 -9508 386 -9212
rect -307 -9560 15 -9559
rect -307 -9880 -306 -9560
rect 14 -9880 15 -9560
rect -307 -9881 15 -9880
rect -198 -10279 -94 -9881
rect 282 -9932 302 -9508
rect 366 -9932 386 -9508
rect 282 -10228 386 -9932
rect -307 -10280 15 -10279
rect -307 -10600 -306 -10280
rect 14 -10600 15 -10280
rect -307 -10601 15 -10600
rect -198 -10999 -94 -10601
rect 282 -10652 302 -10228
rect 366 -10652 386 -10228
rect 282 -10948 386 -10652
rect -307 -11000 15 -10999
rect -307 -11320 -306 -11000
rect 14 -11320 15 -11000
rect -307 -11321 15 -11320
rect -198 -11719 -94 -11321
rect 282 -11372 302 -10948
rect 366 -11372 386 -10948
rect 282 -11668 386 -11372
rect -307 -11720 15 -11719
rect -307 -12040 -306 -11720
rect 14 -12040 15 -11720
rect -307 -12041 15 -12040
rect -198 -12439 -94 -12041
rect 282 -12092 302 -11668
rect 366 -12092 386 -11668
rect 282 -12388 386 -12092
rect -307 -12440 15 -12439
rect -307 -12760 -306 -12440
rect 14 -12760 15 -12440
rect -307 -12761 15 -12760
rect -198 -13159 -94 -12761
rect 282 -12812 302 -12388
rect 366 -12812 386 -12388
rect 282 -13108 386 -12812
rect -307 -13160 15 -13159
rect -307 -13480 -306 -13160
rect 14 -13480 15 -13160
rect -307 -13481 15 -13480
rect -198 -13879 -94 -13481
rect 282 -13532 302 -13108
rect 366 -13532 386 -13108
rect 282 -13828 386 -13532
rect -307 -13880 15 -13879
rect -307 -14200 -306 -13880
rect 14 -14200 15 -13880
rect -307 -14201 15 -14200
rect -198 -14599 -94 -14201
rect 282 -14252 302 -13828
rect 366 -14252 386 -13828
rect 282 -14548 386 -14252
rect -307 -14600 15 -14599
rect -307 -14920 -306 -14600
rect 14 -14920 15 -14600
rect -307 -14921 15 -14920
rect -198 -15319 -94 -14921
rect 282 -14972 302 -14548
rect 366 -14972 386 -14548
rect 282 -15268 386 -14972
rect -307 -15320 15 -15319
rect -307 -15640 -306 -15320
rect 14 -15640 15 -15320
rect -307 -15641 15 -15640
rect -198 -16039 -94 -15641
rect 282 -15692 302 -15268
rect 366 -15692 386 -15268
rect 282 -15988 386 -15692
rect -307 -16040 15 -16039
rect -307 -16360 -306 -16040
rect 14 -16360 15 -16040
rect -307 -16361 15 -16360
rect -198 -16759 -94 -16361
rect 282 -16412 302 -15988
rect 366 -16412 386 -15988
rect 282 -16708 386 -16412
rect -307 -16760 15 -16759
rect -307 -17080 -306 -16760
rect 14 -17080 15 -16760
rect -307 -17081 15 -17080
rect -198 -17479 -94 -17081
rect 282 -17132 302 -16708
rect 366 -17132 386 -16708
rect 282 -17428 386 -17132
rect -307 -17480 15 -17479
rect -307 -17800 -306 -17480
rect 14 -17800 15 -17480
rect -307 -17801 15 -17800
rect -198 -18199 -94 -17801
rect 282 -17852 302 -17428
rect 366 -17852 386 -17428
rect 282 -18148 386 -17852
rect -307 -18200 15 -18199
rect -307 -18520 -306 -18200
rect 14 -18520 15 -18200
rect -307 -18521 15 -18520
rect -198 -18919 -94 -18521
rect 282 -18572 302 -18148
rect 366 -18572 386 -18148
rect 282 -18868 386 -18572
rect -307 -18920 15 -18919
rect -307 -19240 -306 -18920
rect 14 -19240 15 -18920
rect -307 -19241 15 -19240
rect -198 -19639 -94 -19241
rect 282 -19292 302 -18868
rect 366 -19292 386 -18868
rect 282 -19588 386 -19292
rect -307 -19640 15 -19639
rect -307 -19960 -306 -19640
rect 14 -19960 15 -19640
rect -307 -19961 15 -19960
rect -198 -20359 -94 -19961
rect 282 -20012 302 -19588
rect 366 -20012 386 -19588
rect 282 -20308 386 -20012
rect -307 -20360 15 -20359
rect -307 -20680 -306 -20360
rect 14 -20680 15 -20360
rect -307 -20681 15 -20680
rect -198 -21079 -94 -20681
rect 282 -20732 302 -20308
rect 366 -20732 386 -20308
rect 282 -21028 386 -20732
rect -307 -21080 15 -21079
rect -307 -21400 -306 -21080
rect 14 -21400 15 -21080
rect -307 -21401 15 -21400
rect -198 -21799 -94 -21401
rect 282 -21452 302 -21028
rect 366 -21452 386 -21028
rect 282 -21748 386 -21452
rect -307 -21800 15 -21799
rect -307 -22120 -306 -21800
rect 14 -22120 15 -21800
rect -307 -22121 15 -22120
rect -198 -22519 -94 -22121
rect 282 -22172 302 -21748
rect 366 -22172 386 -21748
rect 282 -22468 386 -22172
rect -307 -22520 15 -22519
rect -307 -22840 -306 -22520
rect 14 -22840 15 -22520
rect -307 -22841 15 -22840
rect -198 -23239 -94 -22841
rect 282 -22892 302 -22468
rect 366 -22892 386 -22468
rect 282 -23188 386 -22892
rect -307 -23240 15 -23239
rect -307 -23560 -306 -23240
rect 14 -23560 15 -23240
rect -307 -23561 15 -23560
rect -198 -23959 -94 -23561
rect 282 -23612 302 -23188
rect 366 -23612 386 -23188
rect 282 -23908 386 -23612
rect -307 -23960 15 -23959
rect -307 -24280 -306 -23960
rect 14 -24280 15 -23960
rect -307 -24281 15 -24280
rect -198 -24679 -94 -24281
rect 282 -24332 302 -23908
rect 366 -24332 386 -23908
rect 282 -24628 386 -24332
rect -307 -24680 15 -24679
rect -307 -25000 -306 -24680
rect 14 -25000 15 -24680
rect -307 -25001 15 -25000
rect -198 -25399 -94 -25001
rect 282 -25052 302 -24628
rect 366 -25052 386 -24628
rect 282 -25348 386 -25052
rect -307 -25400 15 -25399
rect -307 -25720 -306 -25400
rect 14 -25720 15 -25400
rect -307 -25721 15 -25720
rect -198 -26119 -94 -25721
rect 282 -25772 302 -25348
rect 366 -25772 386 -25348
rect 282 -26068 386 -25772
rect -307 -26120 15 -26119
rect -307 -26440 -306 -26120
rect 14 -26440 15 -26120
rect -307 -26441 15 -26440
rect -198 -26839 -94 -26441
rect 282 -26492 302 -26068
rect 366 -26492 386 -26068
rect 282 -26788 386 -26492
rect -307 -26840 15 -26839
rect -307 -27160 -306 -26840
rect 14 -27160 15 -26840
rect -307 -27161 15 -27160
rect -198 -27559 -94 -27161
rect 282 -27212 302 -26788
rect 366 -27212 386 -26788
rect 282 -27508 386 -27212
rect -307 -27560 15 -27559
rect -307 -27880 -306 -27560
rect 14 -27880 15 -27560
rect -307 -27881 15 -27880
rect -198 -28279 -94 -27881
rect 282 -27932 302 -27508
rect 366 -27932 386 -27508
rect 282 -28228 386 -27932
rect -307 -28280 15 -28279
rect -307 -28600 -306 -28280
rect 14 -28600 15 -28280
rect -307 -28601 15 -28600
rect -198 -28999 -94 -28601
rect 282 -28652 302 -28228
rect 366 -28652 386 -28228
rect 282 -28948 386 -28652
rect -307 -29000 15 -28999
rect -307 -29320 -306 -29000
rect 14 -29320 15 -29000
rect -307 -29321 15 -29320
rect -198 -29719 -94 -29321
rect 282 -29372 302 -28948
rect 366 -29372 386 -28948
rect 282 -29668 386 -29372
rect -307 -29720 15 -29719
rect -307 -30040 -306 -29720
rect 14 -30040 15 -29720
rect -307 -30041 15 -30040
rect -198 -30439 -94 -30041
rect 282 -30092 302 -29668
rect 366 -30092 386 -29668
rect 282 -30388 386 -30092
rect -307 -30440 15 -30439
rect -307 -30760 -306 -30440
rect 14 -30760 15 -30440
rect -307 -30761 15 -30760
rect -198 -31159 -94 -30761
rect 282 -30812 302 -30388
rect 366 -30812 386 -30388
rect 282 -31108 386 -30812
rect -307 -31160 15 -31159
rect -307 -31480 -306 -31160
rect 14 -31480 15 -31160
rect -307 -31481 15 -31480
rect -198 -31879 -94 -31481
rect 282 -31532 302 -31108
rect 366 -31532 386 -31108
rect 282 -31828 386 -31532
rect -307 -31880 15 -31879
rect -307 -32200 -306 -31880
rect 14 -32200 15 -31880
rect -307 -32201 15 -32200
rect -198 -32599 -94 -32201
rect 282 -32252 302 -31828
rect 366 -32252 386 -31828
rect 282 -32548 386 -32252
rect -307 -32600 15 -32599
rect -307 -32920 -306 -32600
rect 14 -32920 15 -32600
rect -307 -32921 15 -32920
rect -198 -33319 -94 -32921
rect 282 -32972 302 -32548
rect 366 -32972 386 -32548
rect 282 -33268 386 -32972
rect -307 -33320 15 -33319
rect -307 -33640 -306 -33320
rect 14 -33640 15 -33320
rect -307 -33641 15 -33640
rect -198 -34039 -94 -33641
rect 282 -33692 302 -33268
rect 366 -33692 386 -33268
rect 282 -33988 386 -33692
rect -307 -34040 15 -34039
rect -307 -34360 -306 -34040
rect 14 -34360 15 -34040
rect -307 -34361 15 -34360
rect -198 -34759 -94 -34361
rect 282 -34412 302 -33988
rect 366 -34412 386 -33988
rect 282 -34708 386 -34412
rect -307 -34760 15 -34759
rect -307 -35080 -306 -34760
rect 14 -35080 15 -34760
rect -307 -35081 15 -35080
rect -198 -35479 -94 -35081
rect 282 -35132 302 -34708
rect 366 -35132 386 -34708
rect 282 -35428 386 -35132
rect -307 -35480 15 -35479
rect -307 -35800 -306 -35480
rect 14 -35800 15 -35480
rect -307 -35801 15 -35800
rect -198 -36199 -94 -35801
rect 282 -35852 302 -35428
rect 366 -35852 386 -35428
rect 282 -36148 386 -35852
rect -307 -36200 15 -36199
rect -307 -36520 -306 -36200
rect 14 -36520 15 -36200
rect -307 -36521 15 -36520
rect -198 -36919 -94 -36521
rect 282 -36572 302 -36148
rect 366 -36572 386 -36148
rect 282 -36868 386 -36572
rect -307 -36920 15 -36919
rect -307 -37240 -306 -36920
rect 14 -37240 15 -36920
rect -307 -37241 15 -37240
rect -198 -37639 -94 -37241
rect 282 -37292 302 -36868
rect 366 -37292 386 -36868
rect 282 -37588 386 -37292
rect -307 -37640 15 -37639
rect -307 -37960 -306 -37640
rect 14 -37960 15 -37640
rect -307 -37961 15 -37960
rect -198 -38359 -94 -37961
rect 282 -38012 302 -37588
rect 366 -38012 386 -37588
rect 282 -38308 386 -38012
rect -307 -38360 15 -38359
rect -307 -38680 -306 -38360
rect 14 -38680 15 -38360
rect -307 -38681 15 -38680
rect -198 -39079 -94 -38681
rect 282 -38732 302 -38308
rect 366 -38732 386 -38308
rect 282 -39028 386 -38732
rect -307 -39080 15 -39079
rect -307 -39400 -306 -39080
rect 14 -39400 15 -39080
rect -307 -39401 15 -39400
rect -198 -39799 -94 -39401
rect 282 -39452 302 -39028
rect 366 -39452 386 -39028
rect 282 -39748 386 -39452
rect -307 -39800 15 -39799
rect -307 -40120 -306 -39800
rect 14 -40120 15 -39800
rect -307 -40121 15 -40120
rect -198 -40519 -94 -40121
rect 282 -40172 302 -39748
rect 366 -40172 386 -39748
rect 282 -40468 386 -40172
rect -307 -40520 15 -40519
rect -307 -40840 -306 -40520
rect 14 -40840 15 -40520
rect -307 -40841 15 -40840
rect -198 -41239 -94 -40841
rect 282 -40892 302 -40468
rect 366 -40892 386 -40468
rect 282 -41188 386 -40892
rect -307 -41240 15 -41239
rect -307 -41560 -306 -41240
rect 14 -41560 15 -41240
rect -307 -41561 15 -41560
rect -198 -41959 -94 -41561
rect 282 -41612 302 -41188
rect 366 -41612 386 -41188
rect 282 -41908 386 -41612
rect -307 -41960 15 -41959
rect -307 -42280 -306 -41960
rect 14 -42280 15 -41960
rect -307 -42281 15 -42280
rect -198 -42679 -94 -42281
rect 282 -42332 302 -41908
rect 366 -42332 386 -41908
rect 282 -42628 386 -42332
rect -307 -42680 15 -42679
rect -307 -43000 -306 -42680
rect 14 -43000 15 -42680
rect -307 -43001 15 -43000
rect -198 -43399 -94 -43001
rect 282 -43052 302 -42628
rect 366 -43052 386 -42628
rect 282 -43348 386 -43052
rect -307 -43400 15 -43399
rect -307 -43720 -306 -43400
rect 14 -43720 15 -43400
rect -307 -43721 15 -43720
rect -198 -44119 -94 -43721
rect 282 -43772 302 -43348
rect 366 -43772 386 -43348
rect 282 -44068 386 -43772
rect -307 -44120 15 -44119
rect -307 -44440 -306 -44120
rect 14 -44440 15 -44120
rect -307 -44441 15 -44440
rect -198 -44839 -94 -44441
rect 282 -44492 302 -44068
rect 366 -44492 386 -44068
rect 282 -44788 386 -44492
rect -307 -44840 15 -44839
rect -307 -45160 -306 -44840
rect 14 -45160 15 -44840
rect -307 -45161 15 -45160
rect -198 -45559 -94 -45161
rect 282 -45212 302 -44788
rect 366 -45212 386 -44788
rect 282 -45508 386 -45212
rect -307 -45560 15 -45559
rect -307 -45880 -306 -45560
rect 14 -45880 15 -45560
rect -307 -45881 15 -45880
rect -198 -46080 -94 -45881
rect 282 -45932 302 -45508
rect 366 -45932 386 -45508
rect 282 -46080 386 -45932
<< properties >>
string FIXED_BBOX -386 45480 94 45960
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.0 l 2.0 val 9.52 carea 2.00 cperi 0.19 nx 1 ny 128 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
