magic
tech sky130A
timestamp 1730907816
<< pwell >>
rect -123 -505 123 505
<< nmos >>
rect -25 -400 25 400
<< ndiff >>
rect -54 394 -25 400
rect -54 -394 -48 394
rect -31 -394 -25 394
rect -54 -400 -25 -394
rect 25 394 54 400
rect 25 -394 31 394
rect 48 -394 54 394
rect 25 -400 54 -394
<< ndiffc >>
rect -48 -394 -31 394
rect 31 -394 48 394
<< psubdiff >>
rect -105 470 -57 487
rect 57 470 105 487
rect -105 439 -88 470
rect 88 439 105 470
rect -105 -470 -88 -439
rect 88 -470 105 -439
rect -105 -487 -57 -470
rect 57 -487 105 -470
<< psubdiffcont >>
rect -57 470 57 487
rect -105 -439 -88 439
rect 88 -439 105 439
rect -57 -487 57 -470
<< poly >>
rect -25 436 25 444
rect -25 419 -17 436
rect 17 419 25 436
rect -25 400 25 419
rect -25 -419 25 -400
rect -25 -436 -17 -419
rect 17 -436 25 -419
rect -25 -444 25 -436
<< polycont >>
rect -17 419 17 436
rect -17 -436 17 -419
<< locali >>
rect -105 470 -57 487
rect 57 470 105 487
rect -105 439 -88 470
rect 88 439 105 470
rect -25 419 -17 436
rect 17 419 25 436
rect -48 394 -31 402
rect -48 -402 -31 -394
rect 31 394 48 402
rect 31 -402 48 -394
rect -25 -436 -17 -419
rect 17 -436 25 -419
rect -105 -470 -88 -439
rect 88 -470 105 -439
rect -105 -487 -57 -470
rect 57 -487 105 -470
<< viali >>
rect -17 419 17 436
rect -48 -394 -31 394
rect 31 -394 48 394
rect -17 -436 17 -419
<< metal1 >>
rect -23 436 23 439
rect -23 419 -17 436
rect 17 419 23 436
rect -23 416 23 419
rect -51 394 -28 400
rect -51 -394 -48 394
rect -31 -394 -28 394
rect -51 -400 -28 -394
rect 28 394 51 400
rect 28 -394 31 394
rect 48 -394 51 394
rect 28 -400 51 -394
rect -23 -419 23 -416
rect -23 -436 -17 -419
rect 17 -436 23 -419
rect -23 -439 23 -436
<< properties >>
string FIXED_BBOX -96 -478 96 478
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 8.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
