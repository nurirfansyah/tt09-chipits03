magic
tech sky130A
magscale 1 2
timestamp 1729760454
<< metal3 >>
rect -892 1292 -120 1320
rect -892 868 -204 1292
rect -140 868 -120 1292
rect -892 840 -120 868
rect 120 1292 892 1320
rect 120 868 808 1292
rect 872 868 892 1292
rect 120 840 892 868
rect -892 572 -120 600
rect -892 148 -204 572
rect -140 148 -120 572
rect -892 120 -120 148
rect 120 572 892 600
rect 120 148 808 572
rect 872 148 892 572
rect 120 120 892 148
rect -892 -148 -120 -120
rect -892 -572 -204 -148
rect -140 -572 -120 -148
rect -892 -600 -120 -572
rect 120 -148 892 -120
rect 120 -572 808 -148
rect 872 -572 892 -148
rect 120 -600 892 -572
rect -892 -868 -120 -840
rect -892 -1292 -204 -868
rect -140 -1292 -120 -868
rect -892 -1320 -120 -1292
rect 120 -868 892 -840
rect 120 -1292 808 -868
rect 872 -1292 892 -868
rect 120 -1320 892 -1292
<< via3 >>
rect -204 868 -140 1292
rect 808 868 872 1292
rect -204 148 -140 572
rect 808 148 872 572
rect -204 -572 -140 -148
rect 808 -572 872 -148
rect -204 -1292 -140 -868
rect 808 -1292 872 -868
<< mimcap >>
rect -852 1240 -452 1280
rect -852 920 -812 1240
rect -492 920 -452 1240
rect -852 880 -452 920
rect 160 1240 560 1280
rect 160 920 200 1240
rect 520 920 560 1240
rect 160 880 560 920
rect -852 520 -452 560
rect -852 200 -812 520
rect -492 200 -452 520
rect -852 160 -452 200
rect 160 520 560 560
rect 160 200 200 520
rect 520 200 560 520
rect 160 160 560 200
rect -852 -200 -452 -160
rect -852 -520 -812 -200
rect -492 -520 -452 -200
rect -852 -560 -452 -520
rect 160 -200 560 -160
rect 160 -520 200 -200
rect 520 -520 560 -200
rect 160 -560 560 -520
rect -852 -920 -452 -880
rect -852 -1240 -812 -920
rect -492 -1240 -452 -920
rect -852 -1280 -452 -1240
rect 160 -920 560 -880
rect 160 -1240 200 -920
rect 520 -1240 560 -920
rect 160 -1280 560 -1240
<< mimcapcontact >>
rect -812 920 -492 1240
rect 200 920 520 1240
rect -812 200 -492 520
rect 200 200 520 520
rect -812 -520 -492 -200
rect 200 -520 520 -200
rect -812 -1240 -492 -920
rect 200 -1240 520 -920
<< metal4 >>
rect -704 1241 -600 1440
rect -224 1292 -120 1440
rect -813 1240 -491 1241
rect -813 920 -812 1240
rect -492 920 -491 1240
rect -813 919 -491 920
rect -704 521 -600 919
rect -224 868 -204 1292
rect -140 868 -120 1292
rect 308 1241 412 1440
rect 788 1292 892 1440
rect 199 1240 521 1241
rect 199 920 200 1240
rect 520 920 521 1240
rect 199 919 521 920
rect -224 572 -120 868
rect -813 520 -491 521
rect -813 200 -812 520
rect -492 200 -491 520
rect -813 199 -491 200
rect -704 -199 -600 199
rect -224 148 -204 572
rect -140 148 -120 572
rect 308 521 412 919
rect 788 868 808 1292
rect 872 868 892 1292
rect 788 572 892 868
rect 199 520 521 521
rect 199 200 200 520
rect 520 200 521 520
rect 199 199 521 200
rect -224 -148 -120 148
rect -813 -200 -491 -199
rect -813 -520 -812 -200
rect -492 -520 -491 -200
rect -813 -521 -491 -520
rect -704 -919 -600 -521
rect -224 -572 -204 -148
rect -140 -572 -120 -148
rect 308 -199 412 199
rect 788 148 808 572
rect 872 148 892 572
rect 788 -148 892 148
rect 199 -200 521 -199
rect 199 -520 200 -200
rect 520 -520 521 -200
rect 199 -521 521 -520
rect -224 -868 -120 -572
rect -813 -920 -491 -919
rect -813 -1240 -812 -920
rect -492 -1240 -491 -920
rect -813 -1241 -491 -1240
rect -704 -1440 -600 -1241
rect -224 -1292 -204 -868
rect -140 -1292 -120 -868
rect 308 -919 412 -521
rect 788 -572 808 -148
rect 872 -572 892 -148
rect 788 -868 892 -572
rect 199 -920 521 -919
rect 199 -1240 200 -920
rect 520 -1240 521 -920
rect 199 -1241 521 -1240
rect -224 -1440 -120 -1292
rect 308 -1440 412 -1241
rect 788 -1292 808 -868
rect 872 -1292 892 -868
rect 788 -1440 892 -1292
<< properties >>
string FIXED_BBOX 120 840 600 1320
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 2 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
