magic
tech sky130A
magscale 1 2
timestamp 1727309470
<< metal3 >>
rect -386 812 386 840
rect -386 -812 302 812
rect 366 -812 386 812
rect -386 -840 386 -812
<< via3 >>
rect 302 -812 366 812
<< mimcap >>
rect -346 760 54 800
rect -346 -760 -306 760
rect 14 -760 54 760
rect -346 -800 54 -760
<< mimcapcontact >>
rect -306 -760 14 760
<< metal4 >>
rect 286 812 382 828
rect -307 760 15 761
rect -307 -760 -306 760
rect 14 -760 15 760
rect -307 -761 15 -760
rect 286 -812 302 812
rect 366 -812 382 812
rect 286 -828 382 -812
<< properties >>
string FIXED_BBOX -386 -840 94 840
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.0 l 8.0 val 35.8 carea 2.00 cperi 0.19 class capacitor nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100 mf 1
string sky130_fd_pr__cap_mim_m3_1_RM3YWL parameters
<< end >>
